LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_unsigned.all;

ENTITY decision IS PORT(
     start_pa,clk,rst           :in std_logic;
     iter_max          :in    std_logic_vector(4 downto 0);
     x1            :in std_logic;
     x2            :in std_logic;
     x3            :in std_logic;
     x4            :in std_logic;
     x5            :in std_logic;
     x6            :in std_logic;
     x7            :in std_logic;
     x8            :in std_logic;
     x9            :in std_logic;
     x10            :in std_logic;
     x11            :in std_logic;
     x12            :in std_logic;
     x13            :in std_logic;
     x14            :in std_logic;
     x15            :in std_logic;
     x16            :in std_logic;
     x17            :in std_logic;
     x18            :in std_logic;
     x19            :in std_logic;
     x20            :in std_logic;
     x21            :in std_logic;
     x22            :in std_logic;
     x23            :in std_logic;
     x24            :in std_logic;
     x25            :in std_logic;
     x26            :in std_logic;
     x27            :in std_logic;
     x28            :in std_logic;
     x29            :in std_logic;
     x30            :in std_logic;
     x31            :in std_logic;
     x32            :in std_logic;
     x33            :in std_logic;
     x34            :in std_logic;
     x35            :in std_logic;
     x36            :in std_logic;
     x37            :in std_logic;
     x38            :in std_logic;
     x39            :in std_logic;
     x40            :in std_logic;
     x41            :in std_logic;
     x42            :in std_logic;
     x43            :in std_logic;
     x44            :in std_logic;
     x45            :in std_logic;
     x46            :in std_logic;
     x47            :in std_logic;
     x48            :in std_logic;
     x49            :in std_logic;
     x50            :in std_logic;
     x51            :in std_logic;
     x52            :in std_logic;
     x53            :in std_logic;
     x54            :in std_logic;
     x55            :in std_logic;
     x56            :in std_logic;
     x57            :in std_logic;
     x58            :in std_logic;
     x59            :in std_logic;
     x60            :in std_logic;
     x61            :in std_logic;
     x62            :in std_logic;
     x63            :in std_logic;
     x64            :in std_logic;
     x65            :in std_logic;
     x66            :in std_logic;
     x67            :in std_logic;
     x68            :in std_logic;
     x69            :in std_logic;
     x70            :in std_logic;
     x71            :in std_logic;
     x72            :in std_logic;
     x73            :in std_logic;
     x74            :in std_logic;
     x75            :in std_logic;
     x76            :in std_logic;
     x77            :in std_logic;
     x78            :in std_logic;
     x79            :in std_logic;
     x80            :in std_logic;
     x81            :in std_logic;
     x82            :in std_logic;
     x83            :in std_logic;
     x84            :in std_logic;
     x85            :in std_logic;
     x86            :in std_logic;
     x87            :in std_logic;
     x88            :in std_logic;
     x89            :in std_logic;
     x90            :in std_logic;
     x91            :in std_logic;
     x92            :in std_logic;
     x93            :in std_logic;
     x94            :in std_logic;
     x95            :in std_logic;
     x96            :in std_logic;
     x97            :in std_logic;
     x98            :in std_logic;
     x99            :in std_logic;
     x100            :in std_logic;
     x101            :in std_logic;
     x102            :in std_logic;
     x103            :in std_logic;
     x104            :in std_logic;
     x105            :in std_logic;
     x106            :in std_logic;
     x107            :in std_logic;
     x108            :in std_logic;
     x109            :in std_logic;
     x110            :in std_logic;
     x111            :in std_logic;
     x112            :in std_logic;
     x113            :in std_logic;
     x114            :in std_logic;
     x115            :in std_logic;
     x116            :in std_logic;
     x117            :in std_logic;
     x118            :in std_logic;
     x119            :in std_logic;
     x120            :in std_logic;
     x121            :in std_logic;
     x122            :in std_logic;
     x123            :in std_logic;
     x124            :in std_logic;
     x125            :in std_logic;
     x126            :in std_logic;
     x127            :in std_logic;
     x128            :in std_logic;
     x129            :in std_logic;
     x130            :in std_logic;
     x131            :in std_logic;
     x132            :in std_logic;
     x133            :in std_logic;
     x134            :in std_logic;
     x135            :in std_logic;
     x136            :in std_logic;
     x137            :in std_logic;
     x138            :in std_logic;
     x139            :in std_logic;
     x140            :in std_logic;
     x141            :in std_logic;
     x142            :in std_logic;
     x143            :in std_logic;
     x144            :in std_logic;
     x145            :in std_logic;
     x146            :in std_logic;
     x147            :in std_logic;
     x148            :in std_logic;
     x149            :in std_logic;
     x150            :in std_logic;
     x151            :in std_logic;
     x152            :in std_logic;
     x153            :in std_logic;
     x154            :in std_logic;
     x155            :in std_logic;
     x156            :in std_logic;
     x157            :in std_logic;
     x158            :in std_logic;
     x159            :in std_logic;
     x160            :in std_logic;
     x161            :in std_logic;
     x162            :in std_logic;
     x163            :in std_logic;
     x164            :in std_logic;
     x165            :in std_logic;
     x166            :in std_logic;
     x167            :in std_logic;
     x168            :in std_logic;
     x169            :in std_logic;
     x170            :in std_logic;
     x171            :in std_logic;
     x172            :in std_logic;
     x173            :in std_logic;
     x174            :in std_logic;
     x175            :in std_logic;
     x176            :in std_logic;
     x177            :in std_logic;
     x178            :in std_logic;
     x179            :in std_logic;
     x180            :in std_logic;
     x181            :in std_logic;
     x182            :in std_logic;
     x183            :in std_logic;
     x184            :in std_logic;
     x185            :in std_logic;
     x186            :in std_logic;
     x187            :in std_logic;
     x188            :in std_logic;
     x189            :in std_logic;
     x190            :in std_logic;
     x191            :in std_logic;
     x192            :in std_logic;
     x193            :in std_logic;
     x194            :in std_logic;
     x195            :in std_logic;
     x196            :in std_logic;
     x197            :in std_logic;
     x198            :in std_logic;
     x199            :in std_logic;
     x200            :in std_logic;
     x201            :in std_logic;
     x202            :in std_logic;
     x203            :in std_logic;
     x204            :in std_logic;
     x205            :in std_logic;
     x206            :in std_logic;
     x207            :in std_logic;
     x208            :in std_logic;
     x209            :in std_logic;
     x210            :in std_logic;
     x211            :in std_logic;
     x212            :in std_logic;
     x213            :in std_logic;
     x214            :in std_logic;
     x215            :in std_logic;
     x216            :in std_logic;
     x217            :in std_logic;
     x218            :in std_logic;
     x219            :in std_logic;
     x220            :in std_logic;
     x221            :in std_logic;
     x222            :in std_logic;
     x223            :in std_logic;
     x224            :in std_logic;
     x225            :in std_logic;
     x226            :in std_logic;
     x227            :in std_logic;
     x228            :in std_logic;
     x229            :in std_logic;
     x230            :in std_logic;
     x231            :in std_logic;
     x232            :in std_logic;
     x233            :in std_logic;
     x234            :in std_logic;
     x235            :in std_logic;
     x236            :in std_logic;
     x237            :in std_logic;
     x238            :in std_logic;
     x239            :in std_logic;
     x240            :in std_logic;
     x241            :in std_logic;
     x242            :in std_logic;
     x243            :in std_logic;
     x244            :in std_logic;
     x245            :in std_logic;
     x246            :in std_logic;
     x247            :in std_logic;
     x248            :in std_logic;
     x249            :in std_logic;
     x250            :in std_logic;
     x251            :in std_logic;
     x252            :in std_logic;
     x253            :in std_logic;
     x254            :in std_logic;
     x255            :in std_logic;
     x256            :in std_logic;
     x257            :in std_logic;
     x258            :in std_logic;
     x259            :in std_logic;
     x260            :in std_logic;
     x261            :in std_logic;
     x262            :in std_logic;
     x263            :in std_logic;
     x264            :in std_logic;
     x265            :in std_logic;
     x266            :in std_logic;
     x267            :in std_logic;
     x268            :in std_logic;
     x269            :in std_logic;
     x270            :in std_logic;
     x271            :in std_logic;
     x272            :in std_logic;
     x273            :in std_logic;
     x274            :in std_logic;
     x275            :in std_logic;
     x276            :in std_logic;
     x277            :in std_logic;
     x278            :in std_logic;
     x279            :in std_logic;
     x280            :in std_logic;
     x281            :in std_logic;
     x282            :in std_logic;
     x283            :in std_logic;
     x284            :in std_logic;
     x285            :in std_logic;
     x286            :in std_logic;
     x287            :in std_logic;
     x288            :in std_logic;
     x289            :in std_logic;
     x290            :in std_logic;
     x291            :in std_logic;
     x292            :in std_logic;
     x293            :in std_logic;
     x294            :in std_logic;
     x295            :in std_logic;
     x296            :in std_logic;
     x297            :in std_logic;
     x298            :in std_logic;
     x299            :in std_logic;
     x300            :in std_logic;
     x301            :in std_logic;
     x302            :in std_logic;
     x303            :in std_logic;
     x304            :in std_logic;
     x305            :in std_logic;
     x306            :in std_logic;
     x307            :in std_logic;
     x308            :in std_logic;
     x309            :in std_logic;
     x310            :in std_logic;
     x311            :in std_logic;
     x312            :in std_logic;
     x313            :in std_logic;
     x314            :in std_logic;
     x315            :in std_logic;
     x316            :in std_logic;
     x317            :in std_logic;
     x318            :in std_logic;
     x319            :in std_logic;
     x320            :in std_logic;
     x321            :in std_logic;
     x322            :in std_logic;
     x323            :in std_logic;
     x324            :in std_logic;
     x325            :in std_logic;
     x326            :in std_logic;
     x327            :in std_logic;
     x328            :in std_logic;
     x329            :in std_logic;
     x330            :in std_logic;
     x331            :in std_logic;
     x332            :in std_logic;
     x333            :in std_logic;
     x334            :in std_logic;
     x335            :in std_logic;
     x336            :in std_logic;
     x337            :in std_logic;
     x338            :in std_logic;
     x339            :in std_logic;
     x340            :in std_logic;
     x341            :in std_logic;
     x342            :in std_logic;
     x343            :in std_logic;
     x344            :in std_logic;
     x345            :in std_logic;
     x346            :in std_logic;
     x347            :in std_logic;
     x348            :in std_logic;
     x349            :in std_logic;
     x350            :in std_logic;
     x351            :in std_logic;
     x352            :in std_logic;
     x353            :in std_logic;
     x354            :in std_logic;
     x355            :in std_logic;
     x356            :in std_logic;
     x357            :in std_logic;
     x358            :in std_logic;
     x359            :in std_logic;
     x360            :in std_logic;
     x361            :in std_logic;
     x362            :in std_logic;
     x363            :in std_logic;
     x364            :in std_logic;
     x365            :in std_logic;
     x366            :in std_logic;
     x367            :in std_logic;
     x368            :in std_logic;
     x369            :in std_logic;
     x370            :in std_logic;
     x371            :in std_logic;
     x372            :in std_logic;
     x373            :in std_logic;
     x374            :in std_logic;
     x375            :in std_logic;
     x376            :in std_logic;
     x377            :in std_logic;
     x378            :in std_logic;
     x379            :in std_logic;
     x380            :in std_logic;
     x381            :in std_logic;
     x382            :in std_logic;
     x383            :in std_logic;
     x384            :in std_logic;
     x385            :in std_logic;
     x386            :in std_logic;
     x387            :in std_logic;
     x388            :in std_logic;
     x389            :in std_logic;
     x390            :in std_logic;
     x391            :in std_logic;
     x392            :in std_logic;
     x393            :in std_logic;
     x394            :in std_logic;
     x395            :in std_logic;
     x396            :in std_logic;
     x397            :in std_logic;
     x398            :in std_logic;
     x399            :in std_logic;
     x400            :in std_logic;
     x401            :in std_logic;
     x402            :in std_logic;
     x403            :in std_logic;
     x404            :in std_logic;
     x405            :in std_logic;
     x406            :in std_logic;
     x407            :in std_logic;
     x408            :in std_logic;
     x409            :in std_logic;
     x410            :in std_logic;
     x411            :in std_logic;
     x412            :in std_logic;
     x413            :in std_logic;
     x414            :in std_logic;
     x415            :in std_logic;
     x416            :in std_logic;
     x417            :in std_logic;
     x418            :in std_logic;
     x419            :in std_logic;
     x420            :in std_logic;
     x421            :in std_logic;
     x422            :in std_logic;
     x423            :in std_logic;
     x424            :in std_logic;
     x425            :in std_logic;
     x426            :in std_logic;
     x427            :in std_logic;
     x428            :in std_logic;
     x429            :in std_logic;
     x430            :in std_logic;
     x431            :in std_logic;
     x432            :in std_logic;
     x433            :in std_logic;
     x434            :in std_logic;
     x435            :in std_logic;
     x436            :in std_logic;
     x437            :in std_logic;
     x438            :in std_logic;
     x439            :in std_logic;
     x440            :in std_logic;
     x441            :in std_logic;
     x442            :in std_logic;
     x443            :in std_logic;
     x444            :in std_logic;
     x445            :in std_logic;
     x446            :in std_logic;
     x447            :in std_logic;
     x448            :in std_logic;
     x449            :in std_logic;
     x450            :in std_logic;
     x451            :in std_logic;
     x452            :in std_logic;
     x453            :in std_logic;
     x454            :in std_logic;
     x455            :in std_logic;
     x456            :in std_logic;
     x457            :in std_logic;
     x458            :in std_logic;
     x459            :in std_logic;
     x460            :in std_logic;
     x461            :in std_logic;
     x462            :in std_logic;
     x463            :in std_logic;
     x464            :in std_logic;
     x465            :in std_logic;
     x466            :in std_logic;
     x467            :in std_logic;
     x468            :in std_logic;
     x469            :in std_logic;
     x470            :in std_logic;
     x471            :in std_logic;
     x472            :in std_logic;
     x473            :in std_logic;
     x474            :in std_logic;
     x475            :in std_logic;
     x476            :in std_logic;
     x477            :in std_logic;
     x478            :in std_logic;
     x479            :in std_logic;
     x480            :in std_logic;
     x481            :in std_logic;
     x482            :in std_logic;
     x483            :in std_logic;
     x484            :in std_logic;
     x485            :in std_logic;
     x486            :in std_logic;
     x487            :in std_logic;
     x488            :in std_logic;
     x489            :in std_logic;
     x490            :in std_logic;
     x491            :in std_logic;
     x492            :in std_logic;
     x493            :in std_logic;
     x494            :in std_logic;
     x495            :in std_logic;
     x496            :in std_logic;
     x497            :in std_logic;
     x498            :in std_logic;
     x499            :in std_logic;
     x500            :in std_logic;
     x501            :in std_logic;
     x502            :in std_logic;
     x503            :in std_logic;
     x504            :in std_logic;
     x505            :in std_logic;
     x506            :in std_logic;
     x507            :in std_logic;
     x508            :in std_logic;
     x509            :in std_logic;
     x510            :in std_logic;
     x511            :in std_logic;
     x512            :in std_logic;
     x513            :in std_logic;
     x514            :in std_logic;
     x515            :in std_logic;
     x516            :in std_logic;
     x517            :in std_logic;
     x518            :in std_logic;
     x519            :in std_logic;
     x520            :in std_logic;
     x521            :in std_logic;
     x522            :in std_logic;
     x523            :in std_logic;
     x524            :in std_logic;
     x525            :in std_logic;
     x526            :in std_logic;
     x527            :in std_logic;
     x528            :in std_logic;
     x529            :in std_logic;
     x530            :in std_logic;
     x531            :in std_logic;
     x532            :in std_logic;
     x533            :in std_logic;
     x534            :in std_logic;
     x535            :in std_logic;
     x536            :in std_logic;
     x537            :in std_logic;
     x538            :in std_logic;
     x539            :in std_logic;
     x540            :in std_logic;
     x541            :in std_logic;
     x542            :in std_logic;
     x543            :in std_logic;
     x544            :in std_logic;
     x545            :in std_logic;
     x546            :in std_logic;
     x547            :in std_logic;
     x548            :in std_logic;
     x549            :in std_logic;
     x550            :in std_logic;
     x551            :in std_logic;
     x552            :in std_logic;
     x553            :in std_logic;
     x554            :in std_logic;
     x555            :in std_logic;
     x556            :in std_logic;
     x557            :in std_logic;
     x558            :in std_logic;
     x559            :in std_logic;
     x560            :in std_logic;
     x561            :in std_logic;
     x562            :in std_logic;
     x563            :in std_logic;
     x564            :in std_logic;
     x565            :in std_logic;
     x566            :in std_logic;
     x567            :in std_logic;
     x568            :in std_logic;
     x569            :in std_logic;
     x570            :in std_logic;
     x571            :in std_logic;
     x572            :in std_logic;
     x573            :in std_logic;
     x574            :in std_logic;
     x575            :in std_logic;
     x576            :in std_logic;
     x577            :in std_logic;
     x578            :in std_logic;
     x579            :in std_logic;
     x580            :in std_logic;
     x581            :in std_logic;
     x582            :in std_logic;
     x583            :in std_logic;
     x584            :in std_logic;
     x585            :in std_logic;
     x586            :in std_logic;
     x587            :in std_logic;
     x588            :in std_logic;
     x589            :in std_logic;
     x590            :in std_logic;
     x591            :in std_logic;
     x592            :in std_logic;
     x593            :in std_logic;
     x594            :in std_logic;
     x595            :in std_logic;
     x596            :in std_logic;
     x597            :in std_logic;
     x598            :in std_logic;
     x599            :in std_logic;
     x600            :in std_logic;
     x601            :in std_logic;
     x602            :in std_logic;
     x603            :in std_logic;
     x604            :in std_logic;
     x605            :in std_logic;
     x606            :in std_logic;
     x607            :in std_logic;
     x608            :in std_logic;
     x609            :in std_logic;
     x610            :in std_logic;
     x611            :in std_logic;
     x612            :in std_logic;
     x613            :in std_logic;
     x614            :in std_logic;
     x615            :in std_logic;
     x616            :in std_logic;
     x617            :in std_logic;
     x618            :in std_logic;
     x619            :in std_logic;
     x620            :in std_logic;
     x621            :in std_logic;
     x622            :in std_logic;
     x623            :in std_logic;
     x624            :in std_logic;
     x625            :in std_logic;
     x626            :in std_logic;
     x627            :in std_logic;
     x628            :in std_logic;
     x629            :in std_logic;
     x630            :in std_logic;
     x631            :in std_logic;
     x632            :in std_logic;
     x633            :in std_logic;
     x634            :in std_logic;
     x635            :in std_logic;
     x636            :in std_logic;
     x637            :in std_logic;
     x638            :in std_logic;
     x639            :in std_logic;
     x640            :in std_logic;
     x641            :in std_logic;
     x642            :in std_logic;
     x643            :in std_logic;
     x644            :in std_logic;
     x645            :in std_logic;
     x646            :in std_logic;
     x647            :in std_logic;
     x648            :in std_logic;
     x649            :in std_logic;
     x650            :in std_logic;
     x651            :in std_logic;
     x652            :in std_logic;
     x653            :in std_logic;
     x654            :in std_logic;
     x655            :in std_logic;
     x656            :in std_logic;
     x657            :in std_logic;
     x658            :in std_logic;
     x659            :in std_logic;
     x660            :in std_logic;
     x661            :in std_logic;
     x662            :in std_logic;
     x663            :in std_logic;
     x664            :in std_logic;
     x665            :in std_logic;
     x666            :in std_logic;
     x667            :in std_logic;
     x668            :in std_logic;
     x669            :in std_logic;
     x670            :in std_logic;
     x671            :in std_logic;
     x672            :in std_logic;
     x673            :in std_logic;
     x674            :in std_logic;
     x675            :in std_logic;
     x676            :in std_logic;
     x677            :in std_logic;
     x678            :in std_logic;
     x679            :in std_logic;
     x680            :in std_logic;
     x681            :in std_logic;
     x682            :in std_logic;
     x683            :in std_logic;
     x684            :in std_logic;
     x685            :in std_logic;
     x686            :in std_logic;
     x687            :in std_logic;
     x688            :in std_logic;
     x689            :in std_logic;
     x690            :in std_logic;
     x691            :in std_logic;
     x692            :in std_logic;
     x693            :in std_logic;
     x694            :in std_logic;
     x695            :in std_logic;
     x696            :in std_logic;
     x697            :in std_logic;
     x698            :in std_logic;
     x699            :in std_logic;
     x700            :in std_logic;
     x701            :in std_logic;
     x702            :in std_logic;
     x703            :in std_logic;
     x704            :in std_logic;
     x705            :in std_logic;
     x706            :in std_logic;
     x707            :in std_logic;
     x708            :in std_logic;
     x709            :in std_logic;
     x710            :in std_logic;
     x711            :in std_logic;
     x712            :in std_logic;
     x713            :in std_logic;
     x714            :in std_logic;
     x715            :in std_logic;
     x716            :in std_logic;
     x717            :in std_logic;
     x718            :in std_logic;
     x719            :in std_logic;
     x720            :in std_logic;
     x721            :in std_logic;
     x722            :in std_logic;
     x723            :in std_logic;
     x724            :in std_logic;
     x725            :in std_logic;
     x726            :in std_logic;
     x727            :in std_logic;
     x728            :in std_logic;
     x729            :in std_logic;
     x730            :in std_logic;
     x731            :in std_logic;
     x732            :in std_logic;
     x733            :in std_logic;
     x734            :in std_logic;
     x735            :in std_logic;
     x736            :in std_logic;
     x737            :in std_logic;
     x738            :in std_logic;
     x739            :in std_logic;
     x740            :in std_logic;
     x741            :in std_logic;
     x742            :in std_logic;
     x743            :in std_logic;
     x744            :in std_logic;
     x745            :in std_logic;
     x746            :in std_logic;
     x747            :in std_logic;
     x748            :in std_logic;
     x749            :in std_logic;
     x750            :in std_logic;
     x751            :in std_logic;
     x752            :in std_logic;
     x753            :in std_logic;
     x754            :in std_logic;
     x755            :in std_logic;
     x756            :in std_logic;
     x757            :in std_logic;
     x758            :in std_logic;
     x759            :in std_logic;
     x760            :in std_logic;
     x761            :in std_logic;
     x762            :in std_logic;
     x763            :in std_logic;
     x764            :in std_logic;
     x765            :in std_logic;
     x766            :in std_logic;
     x767            :in std_logic;
     x768            :in std_logic;
     x769            :in std_logic;
     x770            :in std_logic;
     x771            :in std_logic;
     x772            :in std_logic;
     x773            :in std_logic;
     x774            :in std_logic;
     x775            :in std_logic;
     x776            :in std_logic;
     x777            :in std_logic;
     x778            :in std_logic;
     x779            :in std_logic;
     x780            :in std_logic;
     x781            :in std_logic;
     x782            :in std_logic;
     x783            :in std_logic;
     x784            :in std_logic;
     x785            :in std_logic;
     x786            :in std_logic;
     x787            :in std_logic;
     x788            :in std_logic;
     x789            :in std_logic;
     x790            :in std_logic;
     x791            :in std_logic;
     x792            :in std_logic;
     x793            :in std_logic;
     x794            :in std_logic;
     x795            :in std_logic;
     x796            :in std_logic;
     x797            :in std_logic;
     x798            :in std_logic;
     x799            :in std_logic;
     x800            :in std_logic;
     x801            :in std_logic;
     x802            :in std_logic;
     x803            :in std_logic;
     x804            :in std_logic;
     x805            :in std_logic;
     x806            :in std_logic;
     x807            :in std_logic;
     x808            :in std_logic;
     x809            :in std_logic;
     x810            :in std_logic;
     x811            :in std_logic;
     x812            :in std_logic;
     x813            :in std_logic;
     x814            :in std_logic;
     x815            :in std_logic;
     x816            :in std_logic;
     x817            :in std_logic;
     x818            :in std_logic;
     x819            :in std_logic;
     x820            :in std_logic;
     x821            :in std_logic;
     x822            :in std_logic;
     x823            :in std_logic;
     x824            :in std_logic;
     x825            :in std_logic;
     x826            :in std_logic;
     x827            :in std_logic;
     x828            :in std_logic;
     x829            :in std_logic;
     x830            :in std_logic;
     x831            :in std_logic;
     x832            :in std_logic;
     x833            :in std_logic;
     x834            :in std_logic;
     x835            :in std_logic;
     x836            :in std_logic;
     x837            :in std_logic;
     x838            :in std_logic;
     x839            :in std_logic;
     x840            :in std_logic;
     x841            :in std_logic;
     x842            :in std_logic;
     x843            :in std_logic;
     x844            :in std_logic;
     x845            :in std_logic;
     x846            :in std_logic;
     x847            :in std_logic;
     x848            :in std_logic;
     x849            :in std_logic;
     x850            :in std_logic;
     x851            :in std_logic;
     x852            :in std_logic;
     x853            :in std_logic;
     x854            :in std_logic;
     x855            :in std_logic;
     x856            :in std_logic;
     x857            :in std_logic;
     x858            :in std_logic;
     x859            :in std_logic;
     x860            :in std_logic;
     x861            :in std_logic;
     x862            :in std_logic;
     x863            :in std_logic;
     x864            :in std_logic;
     x865            :in std_logic;
     x866            :in std_logic;
     x867            :in std_logic;
     x868            :in std_logic;
     x869            :in std_logic;
     x870            :in std_logic;
     x871            :in std_logic;
     x872            :in std_logic;
     x873            :in std_logic;
     x874            :in std_logic;
     x875            :in std_logic;
     x876            :in std_logic;
     x877            :in std_logic;
     x878            :in std_logic;
     x879            :in std_logic;
     x880            :in std_logic;
     x881            :in std_logic;
     x882            :in std_logic;
     x883            :in std_logic;
     x884            :in std_logic;
     x885            :in std_logic;
     x886            :in std_logic;
     x887            :in std_logic;
     x888            :in std_logic;
     x889            :in std_logic;
     x890            :in std_logic;
     x891            :in std_logic;
     x892            :in std_logic;
     x893            :in std_logic;
     x894            :in std_logic;
     x895            :in std_logic;
     x896            :in std_logic;
     x897            :in std_logic;
     x898            :in std_logic;
     x899            :in std_logic;
     x900            :in std_logic;
     x901            :in std_logic;
     x902            :in std_logic;
     x903            :in std_logic;
     x904            :in std_logic;
     x905            :in std_logic;
     x906            :in std_logic;
     x907            :in std_logic;
     x908            :in std_logic;
     x909            :in std_logic;
     x910            :in std_logic;
     x911            :in std_logic;
     x912            :in std_logic;
     x913            :in std_logic;
     x914            :in std_logic;
     x915            :in std_logic;
     x916            :in std_logic;
     x917            :in std_logic;
     x918            :in std_logic;
     x919            :in std_logic;
     x920            :in std_logic;
     x921            :in std_logic;
     x922            :in std_logic;
     x923            :in std_logic;
     x924            :in std_logic;
     x925            :in std_logic;
     x926            :in std_logic;
     x927            :in std_logic;
     x928            :in std_logic;
     x929            :in std_logic;
     x930            :in std_logic;
     x931            :in std_logic;
     x932            :in std_logic;
     x933            :in std_logic;
     x934            :in std_logic;
     x935            :in std_logic;
     x936            :in std_logic;
     x937            :in std_logic;
     x938            :in std_logic;
     x939            :in std_logic;
     x940            :in std_logic;
     x941            :in std_logic;
     x942            :in std_logic;
     x943            :in std_logic;
     x944            :in std_logic;
     x945            :in std_logic;
     x946            :in std_logic;
     x947            :in std_logic;
     x948            :in std_logic;
     x949            :in std_logic;
     x950            :in std_logic;
     x951            :in std_logic;
     x952            :in std_logic;
     x953            :in std_logic;
     x954            :in std_logic;
     x955            :in std_logic;
     x956            :in std_logic;
     x957            :in std_logic;
     x958            :in std_logic;
     x959            :in std_logic;
     x960            :in std_logic;
     x961            :in std_logic;
     x962            :in std_logic;
     x963            :in std_logic;
     x964            :in std_logic;
     x965            :in std_logic;
     x966            :in std_logic;
     x967            :in std_logic;
     x968            :in std_logic;
     x969            :in std_logic;
     x970            :in std_logic;
     x971            :in std_logic;
     x972            :in std_logic;
     x973            :in std_logic;
     x974            :in std_logic;
     x975            :in std_logic;
     x976            :in std_logic;
     x977            :in std_logic;
     x978            :in std_logic;
     x979            :in std_logic;
     x980            :in std_logic;
     x981            :in std_logic;
     x982            :in std_logic;
     x983            :in std_logic;
     x984            :in std_logic;
     x985            :in std_logic;
     x986            :in std_logic;
     x987            :in std_logic;
     x988            :in std_logic;
     x989            :in std_logic;
     x990            :in std_logic;
     x991            :in std_logic;
     x992            :in std_logic;
     x993            :in std_logic;
     x994            :in std_logic;
     x995            :in std_logic;
     x996            :in std_logic;
     x997            :in std_logic;
     x998            :in std_logic;
     x999            :in std_logic;
     x1000            :in std_logic;
     x1001            :in std_logic;
     x1002            :in std_logic;
     x1003            :in std_logic;
     x1004            :in std_logic;
     x1005            :in std_logic;
     x1006            :in std_logic;
     x1007            :in std_logic;
     x1008            :in std_logic;
     x1009            :in std_logic;
     x1010            :in std_logic;
     x1011            :in std_logic;
     x1012            :in std_logic;
     x1013            :in std_logic;
     x1014            :in std_logic;
     x1015            :in std_logic;
     x1016            :in std_logic;
     x1017            :in std_logic;
     x1018            :in std_logic;
     x1019            :in std_logic;
     x1020            :in std_logic;
     x1021            :in std_logic;
     x1022            :in std_logic;
     x1023            :in std_logic;
     x1024            :in std_logic;
     x1025            :in std_logic;
     x1026            :in std_logic;
     x1027            :in std_logic;
     x1028            :in std_logic;
     x1029            :in std_logic;
     x1030            :in std_logic;
     x1031            :in std_logic;
     x1032            :in std_logic;
     x1033            :in std_logic;
     x1034            :in std_logic;
     x1035            :in std_logic;
     x1036            :in std_logic;
     x1037            :in std_logic;
     x1038            :in std_logic;
     x1039            :in std_logic;
     x1040            :in std_logic;
     x1041            :in std_logic;
     x1042            :in std_logic;
     x1043            :in std_logic;
     x1044            :in std_logic;
     x1045            :in std_logic;
     x1046            :in std_logic;
     x1047            :in std_logic;
     x1048            :in std_logic;
     x1049            :in std_logic;
     x1050            :in std_logic;
     x1051            :in std_logic;
     x1052            :in std_logic;
     x1053            :in std_logic;
     x1054            :in std_logic;
     x1055            :in std_logic;
     x1056            :in std_logic;
     x1057            :in std_logic;
     x1058            :in std_logic;
     x1059            :in std_logic;
     x1060            :in std_logic;
     x1061            :in std_logic;
     x1062            :in std_logic;
     x1063            :in std_logic;
     x1064            :in std_logic;
     x1065            :in std_logic;
     x1066            :in std_logic;
     x1067            :in std_logic;
     x1068            :in std_logic;
     x1069            :in std_logic;
     x1070            :in std_logic;
     x1071            :in std_logic;
     x1072            :in std_logic;
     x1073            :in std_logic;
     x1074            :in std_logic;
     x1075            :in std_logic;
     x1076            :in std_logic;
     x1077            :in std_logic;
     x1078            :in std_logic;
     x1079            :in std_logic;
     x1080            :in std_logic;
     x1081            :in std_logic;
     x1082            :in std_logic;
     x1083            :in std_logic;
     x1084            :in std_logic;
     x1085            :in std_logic;
     x1086            :in std_logic;
     x1087            :in std_logic;
     x1088            :in std_logic;
     x1089            :in std_logic;
     x1090            :in std_logic;
     x1091            :in std_logic;
     x1092            :in std_logic;
     x1093            :in std_logic;
     x1094            :in std_logic;
     x1095            :in std_logic;
     x1096            :in std_logic;
     x1097            :in std_logic;
     x1098            :in std_logic;
     x1099            :in std_logic;
     x1100            :in std_logic;
     x1101            :in std_logic;
     x1102            :in std_logic;
     x1103            :in std_logic;
     x1104            :in std_logic;
     x1105            :in std_logic;
     x1106            :in std_logic;
     x1107            :in std_logic;
     x1108            :in std_logic;
     x1109            :in std_logic;
     x1110            :in std_logic;
     x1111            :in std_logic;
     x1112            :in std_logic;
     x1113            :in std_logic;
     x1114            :in std_logic;
     x1115            :in std_logic;
     x1116            :in std_logic;
     x1117            :in std_logic;
     x1118            :in std_logic;
     x1119            :in std_logic;
     x1120            :in std_logic;
     x1121            :in std_logic;
     x1122            :in std_logic;
     x1123            :in std_logic;
     x1124            :in std_logic;
     x1125            :in std_logic;
     x1126            :in std_logic;
     x1127            :in std_logic;
     x1128            :in std_logic;
     x1129            :in std_logic;
     x1130            :in std_logic;
     x1131            :in std_logic;
     x1132            :in std_logic;
     x1133            :in std_logic;
     x1134            :in std_logic;
     x1135            :in std_logic;
     x1136            :in std_logic;
     x1137            :in std_logic;
     x1138            :in std_logic;
     x1139            :in std_logic;
     x1140            :in std_logic;
     x1141            :in std_logic;
     x1142            :in std_logic;
     x1143            :in std_logic;
     x1144            :in std_logic;
     x1145            :in std_logic;
     x1146            :in std_logic;
     x1147            :in std_logic;
     x1148            :in std_logic;
     x1149            :in std_logic;
     x1150            :in std_logic;
     x1151            :in std_logic;
     x1152            :in std_logic;
     x1153            :in std_logic;
     x1154            :in std_logic;
     x1155            :in std_logic;
     x1156            :in std_logic;
     x1157            :in std_logic;
     x1158            :in std_logic;
     x1159            :in std_logic;
     x1160            :in std_logic;
     x1161            :in std_logic;
     x1162            :in std_logic;
     x1163            :in std_logic;
     x1164            :in std_logic;
     x1165            :in std_logic;
     x1166            :in std_logic;
     x1167            :in std_logic;
     x1168            :in std_logic;
     x1169            :in std_logic;
     x1170            :in std_logic;
     x1171            :in std_logic;
     x1172            :in std_logic;
     x1173            :in std_logic;
     x1174            :in std_logic;
     x1175            :in std_logic;
     x1176            :in std_logic;
     x1177            :in std_logic;
     x1178            :in std_logic;
     x1179            :in std_logic;
     x1180            :in std_logic;
     x1181            :in std_logic;
     x1182            :in std_logic;
     x1183            :in std_logic;
     x1184            :in std_logic;
     x1185            :in std_logic;
     x1186            :in std_logic;
     x1187            :in std_logic;
     x1188            :in std_logic;
     x1189            :in std_logic;
     x1190            :in std_logic;
     x1191            :in std_logic;
     x1192            :in std_logic;
     x1193            :in std_logic;
     x1194            :in std_logic;
     x1195            :in std_logic;
     x1196            :in std_logic;
     x1197            :in std_logic;
     x1198            :in std_logic;
     x1199            :in std_logic;
     x1200            :in std_logic;
     x1201            :in std_logic;
     x1202            :in std_logic;
     x1203            :in std_logic;
     x1204            :in std_logic;
     x1205            :in std_logic;
     x1206            :in std_logic;
     x1207            :in std_logic;
     x1208            :in std_logic;
     x1209            :in std_logic;
     x1210            :in std_logic;
     x1211            :in std_logic;
     x1212            :in std_logic;
     x1213            :in std_logic;
     x1214            :in std_logic;
     x1215            :in std_logic;
     x1216            :in std_logic;
     x1217            :in std_logic;
     x1218            :in std_logic;
     x1219            :in std_logic;
     x1220            :in std_logic;
     x1221            :in std_logic;
     x1222            :in std_logic;
     x1223            :in std_logic;
     x1224            :in std_logic;
     x1225            :in std_logic;
     x1226            :in std_logic;
     x1227            :in std_logic;
     x1228            :in std_logic;
     x1229            :in std_logic;
     x1230            :in std_logic;
     x1231            :in std_logic;
     x1232            :in std_logic;
     x1233            :in std_logic;
     x1234            :in std_logic;
     x1235            :in std_logic;
     x1236            :in std_logic;
     x1237            :in std_logic;
     x1238            :in std_logic;
     x1239            :in std_logic;
     x1240            :in std_logic;
     x1241            :in std_logic;
     x1242            :in std_logic;
     x1243            :in std_logic;
     x1244            :in std_logic;
     x1245            :in std_logic;
     x1246            :in std_logic;
     x1247            :in std_logic;
     x1248            :in std_logic;
     x1249            :in std_logic;
     x1250            :in std_logic;
     x1251            :in std_logic;
     x1252            :in std_logic;
     x1253            :in std_logic;
     x1254            :in std_logic;
     x1255            :in std_logic;
     x1256            :in std_logic;
     x1257            :in std_logic;
     x1258            :in std_logic;
     x1259            :in std_logic;
     x1260            :in std_logic;
     x1261            :in std_logic;
     x1262            :in std_logic;
     x1263            :in std_logic;
     x1264            :in std_logic;
     x1265            :in std_logic;
     x1266            :in std_logic;
     x1267            :in std_logic;
     x1268            :in std_logic;
     x1269            :in std_logic;
     x1270            :in std_logic;
     x1271            :in std_logic;
     x1272            :in std_logic;
     x1273            :in std_logic;
     x1274            :in std_logic;
     x1275            :in std_logic;
     x1276            :in std_logic;
     x1277            :in std_logic;
     x1278            :in std_logic;
     x1279            :in std_logic;
     x1280            :in std_logic;
     x1281            :in std_logic;
     x1282            :in std_logic;
     x1283            :in std_logic;
     x1284            :in std_logic;
     x1285            :in std_logic;
     x1286            :in std_logic;
     x1287            :in std_logic;
     x1288            :in std_logic;
     x1289            :in std_logic;
     x1290            :in std_logic;
     x1291            :in std_logic;
     x1292            :in std_logic;
     x1293            :in std_logic;
     x1294            :in std_logic;
     x1295            :in std_logic;
     x1296            :in std_logic;
     x1297            :in std_logic;
     x1298            :in std_logic;
     x1299            :in std_logic;
     x1300            :in std_logic;
     x1301            :in std_logic;
     x1302            :in std_logic;
     x1303            :in std_logic;
     x1304            :in std_logic;
     x1305            :in std_logic;
     x1306            :in std_logic;
     x1307            :in std_logic;
     x1308            :in std_logic;
     x1309            :in std_logic;
     x1310            :in std_logic;
     x1311            :in std_logic;
     x1312            :in std_logic;
     x1313            :in std_logic;
     x1314            :in std_logic;
     x1315            :in std_logic;
     x1316            :in std_logic;
     x1317            :in std_logic;
     x1318            :in std_logic;
     x1319            :in std_logic;
     x1320            :in std_logic;
     x1321            :in std_logic;
     x1322            :in std_logic;
     x1323            :in std_logic;
     x1324            :in std_logic;
     x1325            :in std_logic;
     x1326            :in std_logic;
     x1327            :in std_logic;
     x1328            :in std_logic;
     x1329            :in std_logic;
     x1330            :in std_logic;
     x1331            :in std_logic;
     x1332            :in std_logic;
     x1333            :in std_logic;
     x1334            :in std_logic;
     x1335            :in std_logic;
     x1336            :in std_logic;
     x1337            :in std_logic;
     x1338            :in std_logic;
     x1339            :in std_logic;
     x1340            :in std_logic;
     x1341            :in std_logic;
     x1342            :in std_logic;
     x1343            :in std_logic;
     x1344            :in std_logic;
     x1345            :in std_logic;
     x1346            :in std_logic;
     x1347            :in std_logic;
     x1348            :in std_logic;
     x1349            :in std_logic;
     x1350            :in std_logic;
     x1351            :in std_logic;
     x1352            :in std_logic;
     x1353            :in std_logic;
     x1354            :in std_logic;
     x1355            :in std_logic;
     x1356            :in std_logic;
     x1357            :in std_logic;
     x1358            :in std_logic;
     x1359            :in std_logic;
     x1360            :in std_logic;
     x1361            :in std_logic;
     x1362            :in std_logic;
     x1363            :in std_logic;
     x1364            :in std_logic;
     x1365            :in std_logic;
     x1366            :in std_logic;
     x1367            :in std_logic;
     x1368            :in std_logic;
     x1369            :in std_logic;
     x1370            :in std_logic;
     x1371            :in std_logic;
     x1372            :in std_logic;
     x1373            :in std_logic;
     x1374            :in std_logic;
     x1375            :in std_logic;
     x1376            :in std_logic;
     x1377            :in std_logic;
     x1378            :in std_logic;
     x1379            :in std_logic;
     x1380            :in std_logic;
     x1381            :in std_logic;
     x1382            :in std_logic;
     x1383            :in std_logic;
     x1384            :in std_logic;
     x1385            :in std_logic;
     x1386            :in std_logic;
     x1387            :in std_logic;
     x1388            :in std_logic;
     x1389            :in std_logic;
     x1390            :in std_logic;
     x1391            :in std_logic;
     x1392            :in std_logic;
     x1393            :in std_logic;
     x1394            :in std_logic;
     x1395            :in std_logic;
     x1396            :in std_logic;
     x1397            :in std_logic;
     x1398            :in std_logic;
     x1399            :in std_logic;
     x1400            :in std_logic;
     x1401            :in std_logic;
     x1402            :in std_logic;
     x1403            :in std_logic;
     x1404            :in std_logic;
     x1405            :in std_logic;
     x1406            :in std_logic;
     x1407            :in std_logic;
     x1408            :in std_logic;
     x1409            :in std_logic;
     x1410            :in std_logic;
     x1411            :in std_logic;
     x1412            :in std_logic;
     x1413            :in std_logic;
     x1414            :in std_logic;
     x1415            :in std_logic;
     x1416            :in std_logic;
     x1417            :in std_logic;
     x1418            :in std_logic;
     x1419            :in std_logic;
     x1420            :in std_logic;
     x1421            :in std_logic;
     x1422            :in std_logic;
     x1423            :in std_logic;
     x1424            :in std_logic;
     x1425            :in std_logic;
     x1426            :in std_logic;
     x1427            :in std_logic;
     x1428            :in std_logic;
     x1429            :in std_logic;
     x1430            :in std_logic;
     x1431            :in std_logic;
     x1432            :in std_logic;
     x1433            :in std_logic;
     x1434            :in std_logic;
     x1435            :in std_logic;
     x1436            :in std_logic;
     x1437            :in std_logic;
     x1438            :in std_logic;
     x1439            :in std_logic;
     x1440            :in std_logic;
     x1441            :in std_logic;
     x1442            :in std_logic;
     x1443            :in std_logic;
     x1444            :in std_logic;
     x1445            :in std_logic;
     x1446            :in std_logic;
     x1447            :in std_logic;
     x1448            :in std_logic;
     x1449            :in std_logic;
     x1450            :in std_logic;
     x1451            :in std_logic;
     x1452            :in std_logic;
     x1453            :in std_logic;
     x1454            :in std_logic;
     x1455            :in std_logic;
     x1456            :in std_logic;
     x1457            :in std_logic;
     x1458            :in std_logic;
     x1459            :in std_logic;
     x1460            :in std_logic;
     x1461            :in std_logic;
     x1462            :in std_logic;
     x1463            :in std_logic;
     x1464            :in std_logic;
     x1465            :in std_logic;
     x1466            :in std_logic;
     x1467            :in std_logic;
     x1468            :in std_logic;
     x1469            :in std_logic;
     x1470            :in std_logic;
     x1471            :in std_logic;
     x1472            :in std_logic;
     x1473            :in std_logic;
     x1474            :in std_logic;
     x1475            :in std_logic;
     x1476            :in std_logic;
     x1477            :in std_logic;
     x1478            :in std_logic;
     x1479            :in std_logic;
     x1480            :in std_logic;
     x1481            :in std_logic;
     x1482            :in std_logic;
     x1483            :in std_logic;
     x1484            :in std_logic;
     x1485            :in std_logic;
     x1486            :in std_logic;
     x1487            :in std_logic;
     x1488            :in std_logic;
     x1489            :in std_logic;
     x1490            :in std_logic;
     x1491            :in std_logic;
     x1492            :in std_logic;
     x1493            :in std_logic;
     x1494            :in std_logic;
     x1495            :in std_logic;
     x1496            :in std_logic;
     x1497            :in std_logic;
     x1498            :in std_logic;
     x1499            :in std_logic;
     x1500            :in std_logic;
     x1501            :in std_logic;
     x1502            :in std_logic;
     x1503            :in std_logic;
     x1504            :in std_logic;
     x1505            :in std_logic;
     x1506            :in std_logic;
     x1507            :in std_logic;
     x1508            :in std_logic;
     x1509            :in std_logic;
     x1510            :in std_logic;
     x1511            :in std_logic;
     x1512            :in std_logic;
     x1513            :in std_logic;
     x1514            :in std_logic;
     x1515            :in std_logic;
     x1516            :in std_logic;
     x1517            :in std_logic;
     x1518            :in std_logic;
     x1519            :in std_logic;
     x1520            :in std_logic;
     x1521            :in std_logic;
     x1522            :in std_logic;
     x1523            :in std_logic;
     x1524            :in std_logic;
     x1525            :in std_logic;
     x1526            :in std_logic;
     x1527            :in std_logic;
     x1528            :in std_logic;
     x1529            :in std_logic;
     x1530            :in std_logic;
     x1531            :in std_logic;
     x1532            :in std_logic;
     x1533            :in std_logic;
     x1534            :in std_logic;
     x1535            :in std_logic;
     x1536            :in std_logic;
     x1537            :in std_logic;
     x1538            :in std_logic;
     x1539            :in std_logic;
     x1540            :in std_logic;
     x1541            :in std_logic;
     x1542            :in std_logic;
     x1543            :in std_logic;
     x1544            :in std_logic;
     x1545            :in std_logic;
     x1546            :in std_logic;
     x1547            :in std_logic;
     x1548            :in std_logic;
     x1549            :in std_logic;
     x1550            :in std_logic;
     x1551            :in std_logic;
     x1552            :in std_logic;
     x1553            :in std_logic;
     x1554            :in std_logic;
     x1555            :in std_logic;
     x1556            :in std_logic;
     x1557            :in std_logic;
     x1558            :in std_logic;
     x1559            :in std_logic;
     x1560            :in std_logic;
     x1561            :in std_logic;
     x1562            :in std_logic;
     x1563            :in std_logic;
     x1564            :in std_logic;
     x1565            :in std_logic;
     x1566            :in std_logic;
     x1567            :in std_logic;
     x1568            :in std_logic;
     x1569            :in std_logic;
     x1570            :in std_logic;
     x1571            :in std_logic;
     x1572            :in std_logic;
     x1573            :in std_logic;
     x1574            :in std_logic;
     x1575            :in std_logic;
     x1576            :in std_logic;
     x1577            :in std_logic;
     x1578            :in std_logic;
     x1579            :in std_logic;
     x1580            :in std_logic;
     x1581            :in std_logic;
     x1582            :in std_logic;
     x1583            :in std_logic;
     x1584            :in std_logic;
     x1585            :in std_logic;
     x1586            :in std_logic;
     x1587            :in std_logic;
     x1588            :in std_logic;
     x1589            :in std_logic;
     x1590            :in std_logic;
     x1591            :in std_logic;
     x1592            :in std_logic;
     x1593            :in std_logic;
     x1594            :in std_logic;
     x1595            :in std_logic;
     x1596            :in std_logic;
     x1597            :in std_logic;
     x1598            :in std_logic;
     x1599            :in std_logic;
     x1600            :in std_logic;
     x1601            :in std_logic;
     x1602            :in std_logic;
     x1603            :in std_logic;
     x1604            :in std_logic;
     x1605            :in std_logic;
     x1606            :in std_logic;
     x1607            :in std_logic;
     x1608            :in std_logic;
     x1609            :in std_logic;
     x1610            :in std_logic;
     x1611            :in std_logic;
     x1612            :in std_logic;
     x1613            :in std_logic;
     x1614            :in std_logic;
     x1615            :in std_logic;
     x1616            :in std_logic;
     x1617            :in std_logic;
     x1618            :in std_logic;
     x1619            :in std_logic;
     x1620            :in std_logic;
     x1621            :in std_logic;
     x1622            :in std_logic;
     x1623            :in std_logic;
     x1624            :in std_logic;
     x1625            :in std_logic;
     x1626            :in std_logic;
     x1627            :in std_logic;
     x1628            :in std_logic;
     x1629            :in std_logic;
     x1630            :in std_logic;
     x1631            :in std_logic;
     x1632            :in std_logic;
     x1633            :in std_logic;
     x1634            :in std_logic;
     x1635            :in std_logic;
     x1636            :in std_logic;
     x1637            :in std_logic;
     x1638            :in std_logic;
     x1639            :in std_logic;
     x1640            :in std_logic;
     x1641            :in std_logic;
     x1642            :in std_logic;
     x1643            :in std_logic;
     x1644            :in std_logic;
     x1645            :in std_logic;
     x1646            :in std_logic;
     x1647            :in std_logic;
     x1648            :in std_logic;
     x1649            :in std_logic;
     x1650            :in std_logic;
     x1651            :in std_logic;
     x1652            :in std_logic;
     x1653            :in std_logic;
     x1654            :in std_logic;
     x1655            :in std_logic;
     x1656            :in std_logic;
     x1657            :in std_logic;
     x1658            :in std_logic;
     x1659            :in std_logic;
     x1660            :in std_logic;
     x1661            :in std_logic;
     x1662            :in std_logic;
     x1663            :in std_logic;
     x1664            :in std_logic;
     x1665            :in std_logic;
     x1666            :in std_logic;
     x1667            :in std_logic;
     x1668            :in std_logic;
     x1669            :in std_logic;
     x1670            :in std_logic;
     x1671            :in std_logic;
     x1672            :in std_logic;
     x1673            :in std_logic;
     x1674            :in std_logic;
     x1675            :in std_logic;
     x1676            :in std_logic;
     x1677            :in std_logic;
     x1678            :in std_logic;
     x1679            :in std_logic;
     x1680            :in std_logic;
     x1681            :in std_logic;
     x1682            :in std_logic;
     x1683            :in std_logic;
     x1684            :in std_logic;
     x1685            :in std_logic;
     x1686            :in std_logic;
     x1687            :in std_logic;
     x1688            :in std_logic;
     x1689            :in std_logic;
     x1690            :in std_logic;
     x1691            :in std_logic;
     x1692            :in std_logic;
     x1693            :in std_logic;
     x1694            :in std_logic;
     x1695            :in std_logic;
     x1696            :in std_logic;
     x1697            :in std_logic;
     x1698            :in std_logic;
     x1699            :in std_logic;
     x1700            :in std_logic;
     x1701            :in std_logic;
     x1702            :in std_logic;
     x1703            :in std_logic;
     x1704            :in std_logic;
     x1705            :in std_logic;
     x1706            :in std_logic;
     x1707            :in std_logic;
     x1708            :in std_logic;
     x1709            :in std_logic;
     x1710            :in std_logic;
     x1711            :in std_logic;
     x1712            :in std_logic;
     x1713            :in std_logic;
     x1714            :in std_logic;
     x1715            :in std_logic;
     x1716            :in std_logic;
     x1717            :in std_logic;
     x1718            :in std_logic;
     x1719            :in std_logic;
     x1720            :in std_logic;
     x1721            :in std_logic;
     x1722            :in std_logic;
     x1723            :in std_logic;
     x1724            :in std_logic;
     x1725            :in std_logic;
     x1726            :in std_logic;
     x1727            :in std_logic;
     x1728            :in std_logic;
     x1729            :in std_logic;
     x1730            :in std_logic;
     x1731            :in std_logic;
     x1732            :in std_logic;
     x1733            :in std_logic;
     x1734            :in std_logic;
     x1735            :in std_logic;
     x1736            :in std_logic;
     x1737            :in std_logic;
     x1738            :in std_logic;
     x1739            :in std_logic;
     x1740            :in std_logic;
     x1741            :in std_logic;
     x1742            :in std_logic;
     x1743            :in std_logic;
     x1744            :in std_logic;
     x1745            :in std_logic;
     x1746            :in std_logic;
     x1747            :in std_logic;
     x1748            :in std_logic;
     x1749            :in std_logic;
     x1750            :in std_logic;
     x1751            :in std_logic;
     x1752            :in std_logic;
     x1753            :in std_logic;
     x1754            :in std_logic;
     x1755            :in std_logic;
     x1756            :in std_logic;
     x1757            :in std_logic;
     x1758            :in std_logic;
     x1759            :in std_logic;
     x1760            :in std_logic;
     x1761            :in std_logic;
     x1762            :in std_logic;
     x1763            :in std_logic;
     x1764            :in std_logic;
     x1765            :in std_logic;
     x1766            :in std_logic;
     x1767            :in std_logic;
     x1768            :in std_logic;
     x1769            :in std_logic;
     x1770            :in std_logic;
     x1771            :in std_logic;
     x1772            :in std_logic;
     x1773            :in std_logic;
     x1774            :in std_logic;
     x1775            :in std_logic;
     x1776            :in std_logic;
     x1777            :in std_logic;
     x1778            :in std_logic;
     x1779            :in std_logic;
     x1780            :in std_logic;
     x1781            :in std_logic;
     x1782            :in std_logic;
     x1783            :in std_logic;
     x1784            :in std_logic;
     x1785            :in std_logic;
     x1786            :in std_logic;
     x1787            :in std_logic;
     x1788            :in std_logic;
     x1789            :in std_logic;
     x1790            :in std_logic;
     x1791            :in std_logic;
     x1792            :in std_logic;
     x1793            :in std_logic;
     x1794            :in std_logic;
     x1795            :in std_logic;
     x1796            :in std_logic;
     x1797            :in std_logic;
     x1798            :in std_logic;
     x1799            :in std_logic;
     x1800            :in std_logic;
     x1801            :in std_logic;
     x1802            :in std_logic;
     x1803            :in std_logic;
     x1804            :in std_logic;
     x1805            :in std_logic;
     x1806            :in std_logic;
     x1807            :in std_logic;
     x1808            :in std_logic;
     x1809            :in std_logic;
     x1810            :in std_logic;
     x1811            :in std_logic;
     x1812            :in std_logic;
     x1813            :in std_logic;
     x1814            :in std_logic;
     x1815            :in std_logic;
     x1816            :in std_logic;
     x1817            :in std_logic;
     x1818            :in std_logic;
     x1819            :in std_logic;
     x1820            :in std_logic;
     x1821            :in std_logic;
     x1822            :in std_logic;
     x1823            :in std_logic;
     x1824            :in std_logic;
     x1825            :in std_logic;
     x1826            :in std_logic;
     x1827            :in std_logic;
     x1828            :in std_logic;
     x1829            :in std_logic;
     x1830            :in std_logic;
     x1831            :in std_logic;
     x1832            :in std_logic;
     x1833            :in std_logic;
     x1834            :in std_logic;
     x1835            :in std_logic;
     x1836            :in std_logic;
     x1837            :in std_logic;
     x1838            :in std_logic;
     x1839            :in std_logic;
     x1840            :in std_logic;
     x1841            :in std_logic;
     x1842            :in std_logic;
     x1843            :in std_logic;
     x1844            :in std_logic;
     x1845            :in std_logic;
     x1846            :in std_logic;
     x1847            :in std_logic;
     x1848            :in std_logic;
     x1849            :in std_logic;
     x1850            :in std_logic;
     x1851            :in std_logic;
     x1852            :in std_logic;
     x1853            :in std_logic;
     x1854            :in std_logic;
     x1855            :in std_logic;
     x1856            :in std_logic;
     x1857            :in std_logic;
     x1858            :in std_logic;
     x1859            :in std_logic;
     x1860            :in std_logic;
     x1861            :in std_logic;
     x1862            :in std_logic;
     x1863            :in std_logic;
     x1864            :in std_logic;
     x1865            :in std_logic;
     x1866            :in std_logic;
     x1867            :in std_logic;
     x1868            :in std_logic;
     x1869            :in std_logic;
     x1870            :in std_logic;
     x1871            :in std_logic;
     x1872            :in std_logic;
     x1873            :in std_logic;
     x1874            :in std_logic;
     x1875            :in std_logic;
     x1876            :in std_logic;
     x1877            :in std_logic;
     x1878            :in std_logic;
     x1879            :in std_logic;
     x1880            :in std_logic;
     x1881            :in std_logic;
     x1882            :in std_logic;
     x1883            :in std_logic;
     x1884            :in std_logic;
     x1885            :in std_logic;
     x1886            :in std_logic;
     x1887            :in std_logic;
     x1888            :in std_logic;
     x1889            :in std_logic;
     x1890            :in std_logic;
     x1891            :in std_logic;
     x1892            :in std_logic;
     x1893            :in std_logic;
     x1894            :in std_logic;
     x1895            :in std_logic;
     x1896            :in std_logic;
     x1897            :in std_logic;
     x1898            :in std_logic;
     x1899            :in std_logic;
     x1900            :in std_logic;
     x1901            :in std_logic;
     x1902            :in std_logic;
     x1903            :in std_logic;
     x1904            :in std_logic;
     x1905            :in std_logic;
     x1906            :in std_logic;
     x1907            :in std_logic;
     x1908            :in std_logic;
     x1909            :in std_logic;
     x1910            :in std_logic;
     x1911            :in std_logic;
     x1912            :in std_logic;
     x1913            :in std_logic;
     x1914            :in std_logic;
     x1915            :in std_logic;
     x1916            :in std_logic;
     x1917            :in std_logic;
     x1918            :in std_logic;
     x1919            :in std_logic;
     x1920            :in std_logic;
     x1921            :in std_logic;
     x1922            :in std_logic;
     x1923            :in std_logic;
     x1924            :in std_logic;
     x1925            :in std_logic;
     x1926            :in std_logic;
     x1927            :in std_logic;
     x1928            :in std_logic;
     x1929            :in std_logic;
     x1930            :in std_logic;
     x1931            :in std_logic;
     x1932            :in std_logic;
     x1933            :in std_logic;
     x1934            :in std_logic;
     x1935            :in std_logic;
     x1936            :in std_logic;
     x1937            :in std_logic;
     x1938            :in std_logic;
     x1939            :in std_logic;
     x1940            :in std_logic;
     x1941            :in std_logic;
     x1942            :in std_logic;
     x1943            :in std_logic;
     x1944            :in std_logic;
     x1945            :in std_logic;
     x1946            :in std_logic;
     x1947            :in std_logic;
     x1948            :in std_logic;
     x1949            :in std_logic;
     x1950            :in std_logic;
     x1951            :in std_logic;
     x1952            :in std_logic;
     x1953            :in std_logic;
     x1954            :in std_logic;
     x1955            :in std_logic;
     x1956            :in std_logic;
     x1957            :in std_logic;
     x1958            :in std_logic;
     x1959            :in std_logic;
     x1960            :in std_logic;
     x1961            :in std_logic;
     x1962            :in std_logic;
     x1963            :in std_logic;
     x1964            :in std_logic;
     x1965            :in std_logic;
     x1966            :in std_logic;
     x1967            :in std_logic;
     x1968            :in std_logic;
     x1969            :in std_logic;
     x1970            :in std_logic;
     x1971            :in std_logic;
     x1972            :in std_logic;
     x1973            :in std_logic;
     x1974            :in std_logic;
     x1975            :in std_logic;
     x1976            :in std_logic;
     x1977            :in std_logic;
     x1978            :in std_logic;
     x1979            :in std_logic;
     x1980            :in std_logic;
     x1981            :in std_logic;
     x1982            :in std_logic;
     x1983            :in std_logic;
     x1984            :in std_logic;
     x1985            :in std_logic;
     x1986            :in std_logic;
     x1987            :in std_logic;
     x1988            :in std_logic;
     x1989            :in std_logic;
     x1990            :in std_logic;
     x1991            :in std_logic;
     x1992            :in std_logic;
     x1993            :in std_logic;
     x1994            :in std_logic;
     x1995            :in std_logic;
     x1996            :in std_logic;
     x1997            :in std_logic;
     x1998            :in std_logic;
     x1999            :in std_logic;
     x2000            :in std_logic;
     x2001            :in std_logic;
     x2002            :in std_logic;
     x2003            :in std_logic;
     x2004            :in std_logic;
     x2005            :in std_logic;
     x2006            :in std_logic;
     x2007            :in std_logic;
     x2008            :in std_logic;
     x2009            :in std_logic;
     x2010            :in std_logic;
     x2011            :in std_logic;
     x2012            :in std_logic;
     x2013            :in std_logic;
     x2014            :in std_logic;
     x2015            :in std_logic;
     x2016            :in std_logic;
     x2017            :in std_logic;
     x2018            :in std_logic;
     x2019            :in std_logic;
     x2020            :in std_logic;
     x2021            :in std_logic;
     x2022            :in std_logic;
     x2023            :in std_logic;
     x2024            :in std_logic;
     x2025            :in std_logic;
     x2026            :in std_logic;
     x2027            :in std_logic;
     x2028            :in std_logic;
     x2029            :in std_logic;
     x2030            :in std_logic;
     x2031            :in std_logic;
     x2032            :in std_logic;
     x2033            :in std_logic;
     x2034            :in std_logic;
     x2035            :in std_logic;
     x2036            :in std_logic;
     x2037            :in std_logic;
     x2038            :in std_logic;
     x2039            :in std_logic;
     x2040            :in std_logic;
     x2041            :in std_logic;
     x2042            :in std_logic;
     x2043            :in std_logic;
     x2044            :in std_logic;
     x2045            :in std_logic;
     x2046            :in std_logic;
     x2047            :in std_logic;
     x2048            :in std_logic;
     x2049            :in std_logic;
     x2050            :in std_logic;
     x2051            :in std_logic;
     x2052            :in std_logic;
     x2053            :in std_logic;
     x2054            :in std_logic;
     x2055            :in std_logic;
     x2056            :in std_logic;
     x2057            :in std_logic;
     x2058            :in std_logic;
     x2059            :in std_logic;
     x2060            :in std_logic;
     x2061            :in std_logic;
     x2062            :in std_logic;
     x2063            :in std_logic;
     x2064            :in std_logic;
     x2065            :in std_logic;
     x2066            :in std_logic;
     x2067            :in std_logic;
     x2068            :in std_logic;
     x2069            :in std_logic;
     x2070            :in std_logic;
     x2071            :in std_logic;
     x2072            :in std_logic;
     x2073            :in std_logic;
     x2074            :in std_logic;
     x2075            :in std_logic;
     x2076            :in std_logic;
     x2077            :in std_logic;
     x2078            :in std_logic;
     x2079            :in std_logic;
     x2080            :in std_logic;
     x2081            :in std_logic;
     x2082            :in std_logic;
     x2083            :in std_logic;
     x2084            :in std_logic;
     x2085            :in std_logic;
     x2086            :in std_logic;
     x2087            :in std_logic;
     x2088            :in std_logic;
     x2089            :in std_logic;
     x2090            :in std_logic;
     x2091            :in std_logic;
     x2092            :in std_logic;
     x2093            :in std_logic;
     x2094            :in std_logic;
     x2095            :in std_logic;
     x2096            :in std_logic;
     x2097            :in std_logic;
     x2098            :in std_logic;
     x2099            :in std_logic;
     x2100            :in std_logic;
     x2101            :in std_logic;
     x2102            :in std_logic;
     x2103            :in std_logic;
     x2104            :in std_logic;
     x2105            :in std_logic;
     x2106            :in std_logic;
     x2107            :in std_logic;
     x2108            :in std_logic;
     x2109            :in std_logic;
     x2110            :in std_logic;
     x2111            :in std_logic;
     x2112            :in std_logic;
     x2113            :in std_logic;
     x2114            :in std_logic;
     x2115            :in std_logic;
     x2116            :in std_logic;
     x2117            :in std_logic;
     x2118            :in std_logic;
     x2119            :in std_logic;
     x2120            :in std_logic;
     x2121            :in std_logic;
     x2122            :in std_logic;
     x2123            :in std_logic;
     x2124            :in std_logic;
     x2125            :in std_logic;
     x2126            :in std_logic;
     x2127            :in std_logic;
     x2128            :in std_logic;
     x2129            :in std_logic;
     x2130            :in std_logic;
     x2131            :in std_logic;
     x2132            :in std_logic;
     x2133            :in std_logic;
     x2134            :in std_logic;
     x2135            :in std_logic;
     x2136            :in std_logic;
     x2137            :in std_logic;
     x2138            :in std_logic;
     x2139            :in std_logic;
     x2140            :in std_logic;
     x2141            :in std_logic;
     x2142            :in std_logic;
     x2143            :in std_logic;
     x2144            :in std_logic;
     x2145            :in std_logic;
     x2146            :in std_logic;
     x2147            :in std_logic;
     x2148            :in std_logic;
     x2149            :in std_logic;
     x2150            :in std_logic;
     x2151            :in std_logic;
     x2152            :in std_logic;
     x2153            :in std_logic;
     x2154            :in std_logic;
     x2155            :in std_logic;
     x2156            :in std_logic;
     x2157            :in std_logic;
     x2158            :in std_logic;
     x2159            :in std_logic;
     x2160            :in std_logic;
     x2161            :in std_logic;
     x2162            :in std_logic;
     x2163            :in std_logic;
     x2164            :in std_logic;
     x2165            :in std_logic;
     x2166            :in std_logic;
     x2167            :in std_logic;
     x2168            :in std_logic;
     x2169            :in std_logic;
     x2170            :in std_logic;
     x2171            :in std_logic;
     x2172            :in std_logic;
     x2173            :in std_logic;
     x2174            :in std_logic;
     x2175            :in std_logic;
     x2176            :in std_logic;
     x2177            :in std_logic;
     x2178            :in std_logic;
     x2179            :in std_logic;
     x2180            :in std_logic;
     x2181            :in std_logic;
     x2182            :in std_logic;
     x2183            :in std_logic;
     x2184            :in std_logic;
     x2185            :in std_logic;
     x2186            :in std_logic;
     x2187            :in std_logic;
     x2188            :in std_logic;
     x2189            :in std_logic;
     x2190            :in std_logic;
     x2191            :in std_logic;
     x2192            :in std_logic;
     x2193            :in std_logic;
     x2194            :in std_logic;
     x2195            :in std_logic;
     x2196            :in std_logic;
     x2197            :in std_logic;
     x2198            :in std_logic;
     x2199            :in std_logic;
     x2200            :in std_logic;
     x2201            :in std_logic;
     x2202            :in std_logic;
     x2203            :in std_logic;
     x2204            :in std_logic;
     x2205            :in std_logic;
     x2206            :in std_logic;
     x2207            :in std_logic;
     x2208            :in std_logic;
     x2209            :in std_logic;
     x2210            :in std_logic;
     x2211            :in std_logic;
     x2212            :in std_logic;
     x2213            :in std_logic;
     x2214            :in std_logic;
     x2215            :in std_logic;
     x2216            :in std_logic;
     x2217            :in std_logic;
     x2218            :in std_logic;
     x2219            :in std_logic;
     x2220            :in std_logic;
     x2221            :in std_logic;
     x2222            :in std_logic;
     x2223            :in std_logic;
     x2224            :in std_logic;
     x2225            :in std_logic;
     x2226            :in std_logic;
     x2227            :in std_logic;
     x2228            :in std_logic;
     x2229            :in std_logic;
     x2230            :in std_logic;
     x2231            :in std_logic;
     x2232            :in std_logic;
     x2233            :in std_logic;
     x2234            :in std_logic;
     x2235            :in std_logic;
     x2236            :in std_logic;
     x2237            :in std_logic;
     x2238            :in std_logic;
     x2239            :in std_logic;
     x2240            :in std_logic;
     x2241            :in std_logic;
     x2242            :in std_logic;
     x2243            :in std_logic;
     x2244            :in std_logic;
     x2245            :in std_logic;
     x2246            :in std_logic;
     x2247            :in std_logic;
     x2248            :in std_logic;
     x2249            :in std_logic;
     x2250            :in std_logic;
     x2251            :in std_logic;
     x2252            :in std_logic;
     x2253            :in std_logic;
     x2254            :in std_logic;
     x2255            :in std_logic;
     x2256            :in std_logic;
     x2257            :in std_logic;
     x2258            :in std_logic;
     x2259            :in std_logic;
     x2260            :in std_logic;
     x2261            :in std_logic;
     x2262            :in std_logic;
     x2263            :in std_logic;
     x2264            :in std_logic;
     x2265            :in std_logic;
     x2266            :in std_logic;
     x2267            :in std_logic;
     x2268            :in std_logic;
     x2269            :in std_logic;
     x2270            :in std_logic;
     x2271            :in std_logic;
     x2272            :in std_logic;
     x2273            :in std_logic;
     x2274            :in std_logic;
     x2275            :in std_logic;
     x2276            :in std_logic;
     x2277            :in std_logic;
     x2278            :in std_logic;
     x2279            :in std_logic;
     x2280            :in std_logic;
     x2281            :in std_logic;
     x2282            :in std_logic;
     x2283            :in std_logic;
     x2284            :in std_logic;
     x2285            :in std_logic;
     x2286            :in std_logic;
     x2287            :in std_logic;
     x2288            :in std_logic;
     x2289            :in std_logic;
     x2290            :in std_logic;
     x2291            :in std_logic;
     x2292            :in std_logic;
     x2293            :in std_logic;
     x2294            :in std_logic;
     x2295            :in std_logic;
     x2296            :in std_logic;
     x2297            :in std_logic;
     x2298            :in std_logic;
     x2299            :in std_logic;
     x2300            :in std_logic;
     x2301            :in std_logic;
     x2302            :in std_logic;
     x2303            :in std_logic;
     x2304            :in std_logic;
     nbr_iter       : out std_logic_vector(4 downto 0);
     end_decision   :out std_logic
);
END;

ARCHITECTURE arch_decision OF decision IS

signal count             : unsigned(4 downto 0);
signal itmax             : unsigned(4 downto 0);
signal Par             : std_logic;
signal   a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,a32,a33,a34,a35,a36,a37,a38,a39,a40,a41,a42,a43,a44,a45,a46,a47,a48,a49,a50,a51,a52,a53,a54,a55,a56,a57,a58,a59,a60,a61,a62,a63,a64,a65,a66,a67,a68,a69,a70,a71,a72,a73,a74,a75,a76,a77,a78,a79,a80,a81,a82,a83,a84,a85,a86,a87,a88,a89,a90,a91,a92,a93,a94,a95,a96,a97,a98,a99,a100,a101,a102,a103,a104,a105,a106,a107,a108,a109,a110,a111,a112,a113,a114,a115,a116,a117,a118,a119,a120,a121,a122,a123,a124,a125,a126,a127,a128,a129,a130,a131,a132,a133,a134,a135,a136,a137,a138,a139,a140,a141,a142,a143,a144,a145,a146,a147,a148,a149,a150,a151,a152,a153,a154,a155,a156,a157,a158,a159,a160,a161,a162,a163,a164,a165,a166,a167,a168,a169,a170,a171,a172,a173,a174,a175,a176,a177,a178,a179,a180,a181,a182,a183,a184,a185,a186,a187,a188,a189,a190,a191,a192,a193,a194,a195,a196,a197,a198,a199,a200,a201,a202,a203,a204,a205,a206,a207,a208,a209,a210,a211,a212,a213,a214,a215,a216,a217,a218,a219,a220,a221,a222,a223,a224,a225,a226,a227,a228,a229,a230,a231,a232,a233,a234,a235,a236,a237,a238,a239,a240,a241,a242,a243,a244,a245,a246,a247,a248,a249,a250,a251,a252,a253,a254,a255,a256,a257,a258,a259,a260,a261,a262,a263,a264,a265,a266,a267,a268,a269,a270,a271,a272,a273,a274,a275,a276,a277,a278,a279,a280,a281,a282,a283,a284,a285,a286,a287,a288,a289,a290,a291,a292,a293,a294,a295,a296,a297,a298,a299,a300,a301,a302,a303,a304,a305,a306,a307,a308,a309,a310,a311,a312,a313,a314,a315,a316,a317,a318,a319,a320,a321,a322,a323,a324,a325,a326,a327,a328,a329,a330,a331,a332,a333,a334,a335,a336,a337,a338,a339,a340,a341,a342,a343,a344,a345,a346,a347,a348,a349,a350,a351,a352,a353,a354,a355,a356,a357,a358,a359,a360,a361,a362,a363,a364,a365,a366,a367,a368,a369,a370,a371,a372,a373,a374,a375,a376,a377,a378,a379,a380,a381,a382,a383,a384,a385,a386,a387,a388,a389,a390,a391,a392,a393,a394,a395,a396,a397,a398,a399,a400,a401,a402,a403,a404,a405,a406,a407,a408,a409,a410,a411,a412,a413,a414,a415,a416,a417,a418,a419,a420,a421,a422,a423,a424,a425,a426,a427,a428,a429,a430,a431,a432,a433,a434,a435,a436,a437,a438,a439,a440,a441,a442,a443,a444,a445,a446,a447,a448,a449,a450,a451,a452,a453,a454,a455,a456,a457,a458,a459,a460,a461,a462,a463,a464,a465,a466,a467,a468,a469,a470,a471,a472,a473,a474,a475,a476,a477,a478,a479,a480,a481,a482,a483,a484,a485,a486,a487,a488,a489,a490,a491,a492,a493,a494,a495,a496,a497,a498,a499,a500,a501,a502,a503,a504,a505,a506,a507,a508,a509,a510,a511,a512,a513,a514,a515,a516,a517,a518,a519,a520,a521,a522,a523,a524,a525,a526,a527,a528,a529,a530,a531,a532,a533,a534,a535,a536,a537,a538,a539,a540,a541,a542,a543,a544,a545,a546,a547,a548,a549,a550,a551,a552,a553,a554,a555,a556,a557,a558,a559,a560,a561,a562,a563,a564,a565,a566,a567,a568,a569,a570,a571,a572,a573,a574,a575,a576,a577,a578,a579,a580,a581,a582,a583,a584,a585,a586,a587,a588,a589,a590,a591,a592,a593,a594,a595,a596,a597,a598,a599,a600,a601,a602,a603,a604,a605,a606,a607,a608,a609,a610,a611,a612,a613,a614,a615,a616,a617,a618,a619,a620,a621,a622,a623,a624,a625,a626,a627,a628,a629,a630,a631,a632,a633,a634,a635,a636,a637,a638,a639,a640,a641,a642,a643,a644,a645,a646,a647,a648,a649,a650,a651,a652,a653,a654,a655,a656,a657,a658,a659,a660,a661,a662,a663,a664,a665,a666,a667,a668,a669,a670,a671,a672,a673,a674,a675,a676,a677,a678,a679,a680,a681,a682,a683,a684,a685,a686,a687,a688,a689,a690,a691,a692,a693,a694,a695,a696,a697,a698,a699,a700,a701,a702,a703,a704,a705,a706,a707,a708,a709,a710,a711,a712,a713,a714,a715,a716,a717,a718,a719,a720,a721,a722,a723,a724,a725,a726,a727,a728,a729,a730,a731,a732,a733,a734,a735,a736,a737,a738,a739,a740,a741,a742,a743,a744,a745,a746,a747,a748,a749,a750,a751,a752,a753,a754,a755,a756,a757,a758,a759,a760,a761,a762,a763,a764,a765,a766,a767,a768,a769,a770,a771,a772,a773,a774,a775,a776,a777,a778,a779,a780,a781,a782,a783,a784,a785,a786,a787,a788,a789,a790,a791,a792,a793,a794,a795,a796,a797,a798,a799,a800,a801,a802,a803,a804,a805,a806,a807,a808,a809,a810,a811,a812,a813,a814,a815,a816,a817,a818,a819,a820,a821,a822,a823,a824,a825,a826,a827,a828,a829,a830,a831,a832,a833,a834,a835,a836,a837,a838,a839,a840,a841,a842,a843,a844,a845,a846,a847,a848,a849,a850,a851,a852,a853,a854,a855,a856,a857,a858,a859,a860,a861,a862,a863,a864,a865,a866,a867,a868,a869,a870,a871,a872,a873,a874,a875,a876,a877,a878,a879,a880,a881,a882,a883,a884,a885,a886,a887,a888,a889,a890,a891,a892,a893,a894,a895,a896,a897,a898,a899,a900,a901,a902,a903,a904,a905,a906,a907,a908,a909,a910,a911,a912,a913,a914,a915,a916,a917,a918,a919,a920,a921,a922,a923,a924,a925,a926,a927,a928,a929,a930,a931,a932,a933,a934,a935,a936,a937,a938,a939,a940,a941,a942,a943,a944,a945,a946,a947,a948,a949,a950,a951,a952,a953,a954,a955,a956,a957,a958,a959,a960,a961,a962,a963,a964,a965,a966,a967,a968,a969,a970,a971,a972,a973,a974,a975,a976,a977,a978,a979,a980,a981,a982,a983,a984,a985,a986,a987,a988,a989,a990,a991,a992,a993,a994,a995,a996,a997,a998,a999,a1000,a1001,a1002,a1003,a1004,a1005,a1006,a1007,a1008,a1009,a1010,a1011,a1012,a1013,a1014,a1015,a1016,a1017,a1018,a1019,a1020,a1021,a1022,a1023,a1024,a1025,a1026,a1027,a1028,a1029,a1030,a1031,a1032,a1033,a1034,a1035,a1036,a1037,a1038,a1039,a1040,a1041,a1042,a1043,a1044,a1045,a1046,a1047,a1048,a1049,a1050,a1051,a1052,a1053,a1054,a1055,a1056,a1057,a1058,a1059,a1060,a1061,a1062,a1063,a1064,a1065,a1066,a1067,a1068,a1069,a1070,a1071,a1072,a1073,a1074,a1075,a1076,a1077,a1078,a1079,a1080,a1081,a1082,a1083,a1084,a1085,a1086,a1087,a1088,a1089,a1090,a1091,a1092,a1093,a1094,a1095,a1096,a1097,a1098,a1099,a1100,a1101,a1102,a1103,a1104,a1105,a1106,a1107,a1108,a1109,a1110,a1111,a1112,a1113,a1114,a1115,a1116,a1117,a1118,a1119,a1120,a1121,a1122,a1123,a1124,a1125,a1126,a1127,a1128,a1129,a1130,a1131,a1132,a1133,a1134,a1135,a1136,a1137,a1138,a1139,a1140,a1141,a1142,a1143,a1144,a1145,a1146,a1147,a1148,a1149,a1150,a1151,a1152   :std_logic;

begin

itmax<=unsigned(iter_max);

a1<=x191 xor x266 xor x824 xor x948 xor x1160 xor x1249;
a2<=x192 xor x267 xor x825 xor x949 xor x1161 xor x1250;
a3<=x97 xor x268 xor x826 xor x950 xor x1162 xor x1251;
a4<=x98 xor x269 xor x827 xor x951 xor x1163 xor x1252;
a5<=x99 xor x270 xor x828 xor x952 xor x1164 xor x1253;
a6<=x100 xor x271 xor x829 xor x953 xor x1165 xor x1254;
a7<=x101 xor x272 xor x830 xor x954 xor x1166 xor x1255;
a8<=x102 xor x273 xor x831 xor x955 xor x1167 xor x1256;
a9<=x103 xor x274 xor x832 xor x956 xor x1168 xor x1257;
a10<=x104 xor x275 xor x833 xor x957 xor x1169 xor x1258;
a11<=x105 xor x276 xor x834 xor x958 xor x1170 xor x1259;
a12<=x106 xor x277 xor x835 xor x959 xor x1171 xor x1260;
a13<=x107 xor x278 xor x836 xor x960 xor x1172 xor x1261;
a14<=x108 xor x279 xor x837 xor x865 xor x1173 xor x1262;
a15<=x109 xor x280 xor x838 xor x866 xor x1174 xor x1263;
a16<=x110 xor x281 xor x839 xor x867 xor x1175 xor x1264;
a17<=x111 xor x282 xor x840 xor x868 xor x1176 xor x1265;
a18<=x112 xor x283 xor x841 xor x869 xor x1177 xor x1266;
a19<=x113 xor x284 xor x842 xor x870 xor x1178 xor x1267;
a20<=x114 xor x285 xor x843 xor x871 xor x1179 xor x1268;
a21<=x115 xor x286 xor x844 xor x872 xor x1180 xor x1269;
a22<=x116 xor x287 xor x845 xor x873 xor x1181 xor x1270;
a23<=x117 xor x288 xor x846 xor x874 xor x1182 xor x1271;
a24<=x118 xor x193 xor x847 xor x875 xor x1183 xor x1272;
a25<=x119 xor x194 xor x848 xor x876 xor x1184 xor x1273;
a26<=x120 xor x195 xor x849 xor x877 xor x1185 xor x1274;
a27<=x121 xor x196 xor x850 xor x878 xor x1186 xor x1275;
a28<=x122 xor x197 xor x851 xor x879 xor x1187 xor x1276;
a29<=x123 xor x198 xor x852 xor x880 xor x1188 xor x1277;
a30<=x124 xor x199 xor x853 xor x881 xor x1189 xor x1278;
a31<=x125 xor x200 xor x854 xor x882 xor x1190 xor x1279;
a32<=x126 xor x201 xor x855 xor x883 xor x1191 xor x1280;
a33<=x127 xor x202 xor x856 xor x884 xor x1192 xor x1281;
a34<=x128 xor x203 xor x857 xor x885 xor x1193 xor x1282;
a35<=x129 xor x204 xor x858 xor x886 xor x1194 xor x1283;
a36<=x130 xor x205 xor x859 xor x887 xor x1195 xor x1284;
a37<=x131 xor x206 xor x860 xor x888 xor x1196 xor x1285;
a38<=x132 xor x207 xor x861 xor x889 xor x1197 xor x1286;
a39<=x133 xor x208 xor x862 xor x890 xor x1198 xor x1287;
a40<=x134 xor x209 xor x863 xor x891 xor x1199 xor x1288;
a41<=x135 xor x210 xor x864 xor x892 xor x1200 xor x1289;
a42<=x136 xor x211 xor x769 xor x893 xor x1201 xor x1290;
a43<=x137 xor x212 xor x770 xor x894 xor x1202 xor x1291;
a44<=x138 xor x213 xor x771 xor x895 xor x1203 xor x1292;
a45<=x139 xor x214 xor x772 xor x896 xor x1204 xor x1293;
a46<=x140 xor x215 xor x773 xor x897 xor x1205 xor x1294;
a47<=x141 xor x216 xor x774 xor x898 xor x1206 xor x1295;
a48<=x142 xor x217 xor x775 xor x899 xor x1207 xor x1296;
a49<=x143 xor x218 xor x776 xor x900 xor x1208 xor x1297;
a50<=x144 xor x219 xor x777 xor x901 xor x1209 xor x1298;
a51<=x145 xor x220 xor x778 xor x902 xor x1210 xor x1299;
a52<=x146 xor x221 xor x779 xor x903 xor x1211 xor x1300;
a53<=x147 xor x222 xor x780 xor x904 xor x1212 xor x1301;
a54<=x148 xor x223 xor x781 xor x905 xor x1213 xor x1302;
a55<=x149 xor x224 xor x782 xor x906 xor x1214 xor x1303;
a56<=x150 xor x225 xor x783 xor x907 xor x1215 xor x1304;
a57<=x151 xor x226 xor x784 xor x908 xor x1216 xor x1305;
a58<=x152 xor x227 xor x785 xor x909 xor x1217 xor x1306;
a59<=x153 xor x228 xor x786 xor x910 xor x1218 xor x1307;
a60<=x154 xor x229 xor x787 xor x911 xor x1219 xor x1308;
a61<=x155 xor x230 xor x788 xor x912 xor x1220 xor x1309;
a62<=x156 xor x231 xor x789 xor x913 xor x1221 xor x1310;
a63<=x157 xor x232 xor x790 xor x914 xor x1222 xor x1311;
a64<=x158 xor x233 xor x791 xor x915 xor x1223 xor x1312;
a65<=x159 xor x234 xor x792 xor x916 xor x1224 xor x1313;
a66<=x160 xor x235 xor x793 xor x917 xor x1225 xor x1314;
a67<=x161 xor x236 xor x794 xor x918 xor x1226 xor x1315;
a68<=x162 xor x237 xor x795 xor x919 xor x1227 xor x1316;
a69<=x163 xor x238 xor x796 xor x920 xor x1228 xor x1317;
a70<=x164 xor x239 xor x797 xor x921 xor x1229 xor x1318;
a71<=x165 xor x240 xor x798 xor x922 xor x1230 xor x1319;
a72<=x166 xor x241 xor x799 xor x923 xor x1231 xor x1320;
a73<=x167 xor x242 xor x800 xor x924 xor x1232 xor x1321;
a74<=x168 xor x243 xor x801 xor x925 xor x1233 xor x1322;
a75<=x169 xor x244 xor x802 xor x926 xor x1234 xor x1323;
a76<=x170 xor x245 xor x803 xor x927 xor x1235 xor x1324;
a77<=x171 xor x246 xor x804 xor x928 xor x1236 xor x1325;
a78<=x172 xor x247 xor x805 xor x929 xor x1237 xor x1326;
a79<=x173 xor x248 xor x806 xor x930 xor x1238 xor x1327;
a80<=x174 xor x249 xor x807 xor x931 xor x1239 xor x1328;
a81<=x175 xor x250 xor x808 xor x932 xor x1240 xor x1329;
a82<=x176 xor x251 xor x809 xor x933 xor x1241 xor x1330;
a83<=x177 xor x252 xor x810 xor x934 xor x1242 xor x1331;
a84<=x178 xor x253 xor x811 xor x935 xor x1243 xor x1332;
a85<=x179 xor x254 xor x812 xor x936 xor x1244 xor x1333;
a86<=x180 xor x255 xor x813 xor x937 xor x1245 xor x1334;
a87<=x181 xor x256 xor x814 xor x938 xor x1246 xor x1335;
a88<=x182 xor x257 xor x815 xor x939 xor x1247 xor x1336;
a89<=x183 xor x258 xor x816 xor x940 xor x1248 xor x1337;
a90<=x184 xor x259 xor x817 xor x941 xor x1153 xor x1338;
a91<=x185 xor x260 xor x818 xor x942 xor x1154 xor x1339;
a92<=x186 xor x261 xor x819 xor x943 xor x1155 xor x1340;
a93<=x187 xor x262 xor x820 xor x944 xor x1156 xor x1341;
a94<=x188 xor x263 xor x821 xor x945 xor x1157 xor x1342;
a95<=x189 xor x264 xor x822 xor x946 xor x1158 xor x1343;
a96<=x190 xor x265 xor x823 xor x947 xor x1159 xor x1344;
a97<=x124 xor x503 xor x656 xor x682 xor x1069 xor x1249 xor x1345;
a98<=x125 xor x504 xor x657 xor x683 xor x1070 xor x1250 xor x1346;
a99<=x126 xor x505 xor x658 xor x684 xor x1071 xor x1251 xor x1347;
a100<=x127 xor x506 xor x659 xor x685 xor x1072 xor x1252 xor x1348;
a101<=x128 xor x507 xor x660 xor x686 xor x1073 xor x1253 xor x1349;
a102<=x129 xor x508 xor x661 xor x687 xor x1074 xor x1254 xor x1350;
a103<=x130 xor x509 xor x662 xor x688 xor x1075 xor x1255 xor x1351;
a104<=x131 xor x510 xor x663 xor x689 xor x1076 xor x1256 xor x1352;
a105<=x132 xor x511 xor x664 xor x690 xor x1077 xor x1257 xor x1353;
a106<=x133 xor x512 xor x665 xor x691 xor x1078 xor x1258 xor x1354;
a107<=x134 xor x513 xor x666 xor x692 xor x1079 xor x1259 xor x1355;
a108<=x135 xor x514 xor x667 xor x693 xor x1080 xor x1260 xor x1356;
a109<=x136 xor x515 xor x668 xor x694 xor x1081 xor x1261 xor x1357;
a110<=x137 xor x516 xor x669 xor x695 xor x1082 xor x1262 xor x1358;
a111<=x138 xor x517 xor x670 xor x696 xor x1083 xor x1263 xor x1359;
a112<=x139 xor x518 xor x671 xor x697 xor x1084 xor x1264 xor x1360;
a113<=x140 xor x519 xor x672 xor x698 xor x1085 xor x1265 xor x1361;
a114<=x141 xor x520 xor x577 xor x699 xor x1086 xor x1266 xor x1362;
a115<=x142 xor x521 xor x578 xor x700 xor x1087 xor x1267 xor x1363;
a116<=x143 xor x522 xor x579 xor x701 xor x1088 xor x1268 xor x1364;
a117<=x144 xor x523 xor x580 xor x702 xor x1089 xor x1269 xor x1365;
a118<=x145 xor x524 xor x581 xor x703 xor x1090 xor x1270 xor x1366;
a119<=x146 xor x525 xor x582 xor x704 xor x1091 xor x1271 xor x1367;
a120<=x147 xor x526 xor x583 xor x705 xor x1092 xor x1272 xor x1368;
a121<=x148 xor x527 xor x584 xor x706 xor x1093 xor x1273 xor x1369;
a122<=x149 xor x528 xor x585 xor x707 xor x1094 xor x1274 xor x1370;
a123<=x150 xor x529 xor x586 xor x708 xor x1095 xor x1275 xor x1371;
a124<=x151 xor x530 xor x587 xor x709 xor x1096 xor x1276 xor x1372;
a125<=x152 xor x531 xor x588 xor x710 xor x1097 xor x1277 xor x1373;
a126<=x153 xor x532 xor x589 xor x711 xor x1098 xor x1278 xor x1374;
a127<=x154 xor x533 xor x590 xor x712 xor x1099 xor x1279 xor x1375;
a128<=x155 xor x534 xor x591 xor x713 xor x1100 xor x1280 xor x1376;
a129<=x156 xor x535 xor x592 xor x714 xor x1101 xor x1281 xor x1377;
a130<=x157 xor x536 xor x593 xor x715 xor x1102 xor x1282 xor x1378;
a131<=x158 xor x537 xor x594 xor x716 xor x1103 xor x1283 xor x1379;
a132<=x159 xor x538 xor x595 xor x717 xor x1104 xor x1284 xor x1380;
a133<=x160 xor x539 xor x596 xor x718 xor x1105 xor x1285 xor x1381;
a134<=x161 xor x540 xor x597 xor x719 xor x1106 xor x1286 xor x1382;
a135<=x162 xor x541 xor x598 xor x720 xor x1107 xor x1287 xor x1383;
a136<=x163 xor x542 xor x599 xor x721 xor x1108 xor x1288 xor x1384;
a137<=x164 xor x543 xor x600 xor x722 xor x1109 xor x1289 xor x1385;
a138<=x165 xor x544 xor x601 xor x723 xor x1110 xor x1290 xor x1386;
a139<=x166 xor x545 xor x602 xor x724 xor x1111 xor x1291 xor x1387;
a140<=x167 xor x546 xor x603 xor x725 xor x1112 xor x1292 xor x1388;
a141<=x168 xor x547 xor x604 xor x726 xor x1113 xor x1293 xor x1389;
a142<=x169 xor x548 xor x605 xor x727 xor x1114 xor x1294 xor x1390;
a143<=x170 xor x549 xor x606 xor x728 xor x1115 xor x1295 xor x1391;
a144<=x171 xor x550 xor x607 xor x729 xor x1116 xor x1296 xor x1392;
a145<=x172 xor x551 xor x608 xor x730 xor x1117 xor x1297 xor x1393;
a146<=x173 xor x552 xor x609 xor x731 xor x1118 xor x1298 xor x1394;
a147<=x174 xor x553 xor x610 xor x732 xor x1119 xor x1299 xor x1395;
a148<=x175 xor x554 xor x611 xor x733 xor x1120 xor x1300 xor x1396;
a149<=x176 xor x555 xor x612 xor x734 xor x1121 xor x1301 xor x1397;
a150<=x177 xor x556 xor x613 xor x735 xor x1122 xor x1302 xor x1398;
a151<=x178 xor x557 xor x614 xor x736 xor x1123 xor x1303 xor x1399;
a152<=x179 xor x558 xor x615 xor x737 xor x1124 xor x1304 xor x1400;
a153<=x180 xor x559 xor x616 xor x738 xor x1125 xor x1305 xor x1401;
a154<=x181 xor x560 xor x617 xor x739 xor x1126 xor x1306 xor x1402;
a155<=x182 xor x561 xor x618 xor x740 xor x1127 xor x1307 xor x1403;
a156<=x183 xor x562 xor x619 xor x741 xor x1128 xor x1308 xor x1404;
a157<=x184 xor x563 xor x620 xor x742 xor x1129 xor x1309 xor x1405;
a158<=x185 xor x564 xor x621 xor x743 xor x1130 xor x1310 xor x1406;
a159<=x186 xor x565 xor x622 xor x744 xor x1131 xor x1311 xor x1407;
a160<=x187 xor x566 xor x623 xor x745 xor x1132 xor x1312 xor x1408;
a161<=x188 xor x567 xor x624 xor x746 xor x1133 xor x1313 xor x1409;
a162<=x189 xor x568 xor x625 xor x747 xor x1134 xor x1314 xor x1410;
a163<=x190 xor x569 xor x626 xor x748 xor x1135 xor x1315 xor x1411;
a164<=x191 xor x570 xor x627 xor x749 xor x1136 xor x1316 xor x1412;
a165<=x192 xor x571 xor x628 xor x750 xor x1137 xor x1317 xor x1413;
a166<=x97 xor x572 xor x629 xor x751 xor x1138 xor x1318 xor x1414;
a167<=x98 xor x573 xor x630 xor x752 xor x1139 xor x1319 xor x1415;
a168<=x99 xor x574 xor x631 xor x753 xor x1140 xor x1320 xor x1416;
a169<=x100 xor x575 xor x632 xor x754 xor x1141 xor x1321 xor x1417;
a170<=x101 xor x576 xor x633 xor x755 xor x1142 xor x1322 xor x1418;
a171<=x102 xor x481 xor x634 xor x756 xor x1143 xor x1323 xor x1419;
a172<=x103 xor x482 xor x635 xor x757 xor x1144 xor x1324 xor x1420;
a173<=x104 xor x483 xor x636 xor x758 xor x1145 xor x1325 xor x1421;
a174<=x105 xor x484 xor x637 xor x759 xor x1146 xor x1326 xor x1422;
a175<=x106 xor x485 xor x638 xor x760 xor x1147 xor x1327 xor x1423;
a176<=x107 xor x486 xor x639 xor x761 xor x1148 xor x1328 xor x1424;
a177<=x108 xor x487 xor x640 xor x762 xor x1149 xor x1329 xor x1425;
a178<=x109 xor x488 xor x641 xor x763 xor x1150 xor x1330 xor x1426;
a179<=x110 xor x489 xor x642 xor x764 xor x1151 xor x1331 xor x1427;
a180<=x111 xor x490 xor x643 xor x765 xor x1152 xor x1332 xor x1428;
a181<=x112 xor x491 xor x644 xor x766 xor x1057 xor x1333 xor x1429;
a182<=x113 xor x492 xor x645 xor x767 xor x1058 xor x1334 xor x1430;
a183<=x114 xor x493 xor x646 xor x768 xor x1059 xor x1335 xor x1431;
a184<=x115 xor x494 xor x647 xor x673 xor x1060 xor x1336 xor x1432;
a185<=x116 xor x495 xor x648 xor x674 xor x1061 xor x1337 xor x1433;
a186<=x117 xor x496 xor x649 xor x675 xor x1062 xor x1338 xor x1434;
a187<=x118 xor x497 xor x650 xor x676 xor x1063 xor x1339 xor x1435;
a188<=x119 xor x498 xor x651 xor x677 xor x1064 xor x1340 xor x1436;
a189<=x120 xor x499 xor x652 xor x678 xor x1065 xor x1341 xor x1437;
a190<=x121 xor x500 xor x653 xor x679 xor x1066 xor x1342 xor x1438;
a191<=x122 xor x501 xor x654 xor x680 xor x1067 xor x1343 xor x1439;
a192<=x123 xor x502 xor x655 xor x681 xor x1068 xor x1344 xor x1440;
a193<=x313 xor x407 xor x562 xor x706 xor x1057 xor x1345 xor x1441;
a194<=x314 xor x408 xor x563 xor x707 xor x1058 xor x1346 xor x1442;
a195<=x315 xor x409 xor x564 xor x708 xor x1059 xor x1347 xor x1443;
a196<=x316 xor x410 xor x565 xor x709 xor x1060 xor x1348 xor x1444;
a197<=x317 xor x411 xor x566 xor x710 xor x1061 xor x1349 xor x1445;
a198<=x318 xor x412 xor x567 xor x711 xor x1062 xor x1350 xor x1446;
a199<=x319 xor x413 xor x568 xor x712 xor x1063 xor x1351 xor x1447;
a200<=x320 xor x414 xor x569 xor x713 xor x1064 xor x1352 xor x1448;
a201<=x321 xor x415 xor x570 xor x714 xor x1065 xor x1353 xor x1449;
a202<=x322 xor x416 xor x571 xor x715 xor x1066 xor x1354 xor x1450;
a203<=x323 xor x417 xor x572 xor x716 xor x1067 xor x1355 xor x1451;
a204<=x324 xor x418 xor x573 xor x717 xor x1068 xor x1356 xor x1452;
a205<=x325 xor x419 xor x574 xor x718 xor x1069 xor x1357 xor x1453;
a206<=x326 xor x420 xor x575 xor x719 xor x1070 xor x1358 xor x1454;
a207<=x327 xor x421 xor x576 xor x720 xor x1071 xor x1359 xor x1455;
a208<=x328 xor x422 xor x481 xor x721 xor x1072 xor x1360 xor x1456;
a209<=x329 xor x423 xor x482 xor x722 xor x1073 xor x1361 xor x1457;
a210<=x330 xor x424 xor x483 xor x723 xor x1074 xor x1362 xor x1458;
a211<=x331 xor x425 xor x484 xor x724 xor x1075 xor x1363 xor x1459;
a212<=x332 xor x426 xor x485 xor x725 xor x1076 xor x1364 xor x1460;
a213<=x333 xor x427 xor x486 xor x726 xor x1077 xor x1365 xor x1461;
a214<=x334 xor x428 xor x487 xor x727 xor x1078 xor x1366 xor x1462;
a215<=x335 xor x429 xor x488 xor x728 xor x1079 xor x1367 xor x1463;
a216<=x336 xor x430 xor x489 xor x729 xor x1080 xor x1368 xor x1464;
a217<=x337 xor x431 xor x490 xor x730 xor x1081 xor x1369 xor x1465;
a218<=x338 xor x432 xor x491 xor x731 xor x1082 xor x1370 xor x1466;
a219<=x339 xor x433 xor x492 xor x732 xor x1083 xor x1371 xor x1467;
a220<=x340 xor x434 xor x493 xor x733 xor x1084 xor x1372 xor x1468;
a221<=x341 xor x435 xor x494 xor x734 xor x1085 xor x1373 xor x1469;
a222<=x342 xor x436 xor x495 xor x735 xor x1086 xor x1374 xor x1470;
a223<=x343 xor x437 xor x496 xor x736 xor x1087 xor x1375 xor x1471;
a224<=x344 xor x438 xor x497 xor x737 xor x1088 xor x1376 xor x1472;
a225<=x345 xor x439 xor x498 xor x738 xor x1089 xor x1377 xor x1473;
a226<=x346 xor x440 xor x499 xor x739 xor x1090 xor x1378 xor x1474;
a227<=x347 xor x441 xor x500 xor x740 xor x1091 xor x1379 xor x1475;
a228<=x348 xor x442 xor x501 xor x741 xor x1092 xor x1380 xor x1476;
a229<=x349 xor x443 xor x502 xor x742 xor x1093 xor x1381 xor x1477;
a230<=x350 xor x444 xor x503 xor x743 xor x1094 xor x1382 xor x1478;
a231<=x351 xor x445 xor x504 xor x744 xor x1095 xor x1383 xor x1479;
a232<=x352 xor x446 xor x505 xor x745 xor x1096 xor x1384 xor x1480;
a233<=x353 xor x447 xor x506 xor x746 xor x1097 xor x1385 xor x1481;
a234<=x354 xor x448 xor x507 xor x747 xor x1098 xor x1386 xor x1482;
a235<=x355 xor x449 xor x508 xor x748 xor x1099 xor x1387 xor x1483;
a236<=x356 xor x450 xor x509 xor x749 xor x1100 xor x1388 xor x1484;
a237<=x357 xor x451 xor x510 xor x750 xor x1101 xor x1389 xor x1485;
a238<=x358 xor x452 xor x511 xor x751 xor x1102 xor x1390 xor x1486;
a239<=x359 xor x453 xor x512 xor x752 xor x1103 xor x1391 xor x1487;
a240<=x360 xor x454 xor x513 xor x753 xor x1104 xor x1392 xor x1488;
a241<=x361 xor x455 xor x514 xor x754 xor x1105 xor x1393 xor x1489;
a242<=x362 xor x456 xor x515 xor x755 xor x1106 xor x1394 xor x1490;
a243<=x363 xor x457 xor x516 xor x756 xor x1107 xor x1395 xor x1491;
a244<=x364 xor x458 xor x517 xor x757 xor x1108 xor x1396 xor x1492;
a245<=x365 xor x459 xor x518 xor x758 xor x1109 xor x1397 xor x1493;
a246<=x366 xor x460 xor x519 xor x759 xor x1110 xor x1398 xor x1494;
a247<=x367 xor x461 xor x520 xor x760 xor x1111 xor x1399 xor x1495;
a248<=x368 xor x462 xor x521 xor x761 xor x1112 xor x1400 xor x1496;
a249<=x369 xor x463 xor x522 xor x762 xor x1113 xor x1401 xor x1497;
a250<=x370 xor x464 xor x523 xor x763 xor x1114 xor x1402 xor x1498;
a251<=x371 xor x465 xor x524 xor x764 xor x1115 xor x1403 xor x1499;
a252<=x372 xor x466 xor x525 xor x765 xor x1116 xor x1404 xor x1500;
a253<=x373 xor x467 xor x526 xor x766 xor x1117 xor x1405 xor x1501;
a254<=x374 xor x468 xor x527 xor x767 xor x1118 xor x1406 xor x1502;
a255<=x375 xor x469 xor x528 xor x768 xor x1119 xor x1407 xor x1503;
a256<=x376 xor x470 xor x529 xor x673 xor x1120 xor x1408 xor x1504;
a257<=x377 xor x471 xor x530 xor x674 xor x1121 xor x1409 xor x1505;
a258<=x378 xor x472 xor x531 xor x675 xor x1122 xor x1410 xor x1506;
a259<=x379 xor x473 xor x532 xor x676 xor x1123 xor x1411 xor x1507;
a260<=x380 xor x474 xor x533 xor x677 xor x1124 xor x1412 xor x1508;
a261<=x381 xor x475 xor x534 xor x678 xor x1125 xor x1413 xor x1509;
a262<=x382 xor x476 xor x535 xor x679 xor x1126 xor x1414 xor x1510;
a263<=x383 xor x477 xor x536 xor x680 xor x1127 xor x1415 xor x1511;
a264<=x384 xor x478 xor x537 xor x681 xor x1128 xor x1416 xor x1512;
a265<=x289 xor x479 xor x538 xor x682 xor x1129 xor x1417 xor x1513;
a266<=x290 xor x480 xor x539 xor x683 xor x1130 xor x1418 xor x1514;
a267<=x291 xor x385 xor x540 xor x684 xor x1131 xor x1419 xor x1515;
a268<=x292 xor x386 xor x541 xor x685 xor x1132 xor x1420 xor x1516;
a269<=x293 xor x387 xor x542 xor x686 xor x1133 xor x1421 xor x1517;
a270<=x294 xor x388 xor x543 xor x687 xor x1134 xor x1422 xor x1518;
a271<=x295 xor x389 xor x544 xor x688 xor x1135 xor x1423 xor x1519;
a272<=x296 xor x390 xor x545 xor x689 xor x1136 xor x1424 xor x1520;
a273<=x297 xor x391 xor x546 xor x690 xor x1137 xor x1425 xor x1521;
a274<=x298 xor x392 xor x547 xor x691 xor x1138 xor x1426 xor x1522;
a275<=x299 xor x393 xor x548 xor x692 xor x1139 xor x1427 xor x1523;
a276<=x300 xor x394 xor x549 xor x693 xor x1140 xor x1428 xor x1524;
a277<=x301 xor x395 xor x550 xor x694 xor x1141 xor x1429 xor x1525;
a278<=x302 xor x396 xor x551 xor x695 xor x1142 xor x1430 xor x1526;
a279<=x303 xor x397 xor x552 xor x696 xor x1143 xor x1431 xor x1527;
a280<=x304 xor x398 xor x553 xor x697 xor x1144 xor x1432 xor x1528;
a281<=x305 xor x399 xor x554 xor x698 xor x1145 xor x1433 xor x1529;
a282<=x306 xor x400 xor x555 xor x699 xor x1146 xor x1434 xor x1530;
a283<=x307 xor x401 xor x556 xor x700 xor x1147 xor x1435 xor x1531;
a284<=x308 xor x402 xor x557 xor x701 xor x1148 xor x1436 xor x1532;
a285<=x309 xor x403 xor x558 xor x702 xor x1149 xor x1437 xor x1533;
a286<=x310 xor x404 xor x559 xor x703 xor x1150 xor x1438 xor x1534;
a287<=x311 xor x405 xor x560 xor x704 xor x1151 xor x1439 xor x1535;
a288<=x312 xor x406 xor x561 xor x705 xor x1152 xor x1440 xor x1536;
a289<=x62 xor x240 xor x834 xor x890 xor x1441 xor x1537;
a290<=x63 xor x241 xor x835 xor x891 xor x1442 xor x1538;
a291<=x64 xor x242 xor x836 xor x892 xor x1443 xor x1539;
a292<=x65 xor x243 xor x837 xor x893 xor x1444 xor x1540;
a293<=x66 xor x244 xor x838 xor x894 xor x1445 xor x1541;
a294<=x67 xor x245 xor x839 xor x895 xor x1446 xor x1542;
a295<=x68 xor x246 xor x840 xor x896 xor x1447 xor x1543;
a296<=x69 xor x247 xor x841 xor x897 xor x1448 xor x1544;
a297<=x70 xor x248 xor x842 xor x898 xor x1449 xor x1545;
a298<=x71 xor x249 xor x843 xor x899 xor x1450 xor x1546;
a299<=x72 xor x250 xor x844 xor x900 xor x1451 xor x1547;
a300<=x73 xor x251 xor x845 xor x901 xor x1452 xor x1548;
a301<=x74 xor x252 xor x846 xor x902 xor x1453 xor x1549;
a302<=x75 xor x253 xor x847 xor x903 xor x1454 xor x1550;
a303<=x76 xor x254 xor x848 xor x904 xor x1455 xor x1551;
a304<=x77 xor x255 xor x849 xor x905 xor x1456 xor x1552;
a305<=x78 xor x256 xor x850 xor x906 xor x1457 xor x1553;
a306<=x79 xor x257 xor x851 xor x907 xor x1458 xor x1554;
a307<=x80 xor x258 xor x852 xor x908 xor x1459 xor x1555;
a308<=x81 xor x259 xor x853 xor x909 xor x1460 xor x1556;
a309<=x82 xor x260 xor x854 xor x910 xor x1461 xor x1557;
a310<=x83 xor x261 xor x855 xor x911 xor x1462 xor x1558;
a311<=x84 xor x262 xor x856 xor x912 xor x1463 xor x1559;
a312<=x85 xor x263 xor x857 xor x913 xor x1464 xor x1560;
a313<=x86 xor x264 xor x858 xor x914 xor x1465 xor x1561;
a314<=x87 xor x265 xor x859 xor x915 xor x1466 xor x1562;
a315<=x88 xor x266 xor x860 xor x916 xor x1467 xor x1563;
a316<=x89 xor x267 xor x861 xor x917 xor x1468 xor x1564;
a317<=x90 xor x268 xor x862 xor x918 xor x1469 xor x1565;
a318<=x91 xor x269 xor x863 xor x919 xor x1470 xor x1566;
a319<=x92 xor x270 xor x864 xor x920 xor x1471 xor x1567;
a320<=x93 xor x271 xor x769 xor x921 xor x1472 xor x1568;
a321<=x94 xor x272 xor x770 xor x922 xor x1473 xor x1569;
a322<=x95 xor x273 xor x771 xor x923 xor x1474 xor x1570;
a323<=x96 xor x274 xor x772 xor x924 xor x1475 xor x1571;
a324<=x1 xor x275 xor x773 xor x925 xor x1476 xor x1572;
a325<=x2 xor x276 xor x774 xor x926 xor x1477 xor x1573;
a326<=x3 xor x277 xor x775 xor x927 xor x1478 xor x1574;
a327<=x4 xor x278 xor x776 xor x928 xor x1479 xor x1575;
a328<=x5 xor x279 xor x777 xor x929 xor x1480 xor x1576;
a329<=x6 xor x280 xor x778 xor x930 xor x1481 xor x1577;
a330<=x7 xor x281 xor x779 xor x931 xor x1482 xor x1578;
a331<=x8 xor x282 xor x780 xor x932 xor x1483 xor x1579;
a332<=x9 xor x283 xor x781 xor x933 xor x1484 xor x1580;
a333<=x10 xor x284 xor x782 xor x934 xor x1485 xor x1581;
a334<=x11 xor x285 xor x783 xor x935 xor x1486 xor x1582;
a335<=x12 xor x286 xor x784 xor x936 xor x1487 xor x1583;
a336<=x13 xor x287 xor x785 xor x937 xor x1488 xor x1584;
a337<=x14 xor x288 xor x786 xor x938 xor x1489 xor x1585;
a338<=x15 xor x193 xor x787 xor x939 xor x1490 xor x1586;
a339<=x16 xor x194 xor x788 xor x940 xor x1491 xor x1587;
a340<=x17 xor x195 xor x789 xor x941 xor x1492 xor x1588;
a341<=x18 xor x196 xor x790 xor x942 xor x1493 xor x1589;
a342<=x19 xor x197 xor x791 xor x943 xor x1494 xor x1590;
a343<=x20 xor x198 xor x792 xor x944 xor x1495 xor x1591;
a344<=x21 xor x199 xor x793 xor x945 xor x1496 xor x1592;
a345<=x22 xor x200 xor x794 xor x946 xor x1497 xor x1593;
a346<=x23 xor x201 xor x795 xor x947 xor x1498 xor x1594;
a347<=x24 xor x202 xor x796 xor x948 xor x1499 xor x1595;
a348<=x25 xor x203 xor x797 xor x949 xor x1500 xor x1596;
a349<=x26 xor x204 xor x798 xor x950 xor x1501 xor x1597;
a350<=x27 xor x205 xor x799 xor x951 xor x1502 xor x1598;
a351<=x28 xor x206 xor x800 xor x952 xor x1503 xor x1599;
a352<=x29 xor x207 xor x801 xor x953 xor x1504 xor x1600;
a353<=x30 xor x208 xor x802 xor x954 xor x1505 xor x1601;
a354<=x31 xor x209 xor x803 xor x955 xor x1506 xor x1602;
a355<=x32 xor x210 xor x804 xor x956 xor x1507 xor x1603;
a356<=x33 xor x211 xor x805 xor x957 xor x1508 xor x1604;
a357<=x34 xor x212 xor x806 xor x958 xor x1509 xor x1605;
a358<=x35 xor x213 xor x807 xor x959 xor x1510 xor x1606;
a359<=x36 xor x214 xor x808 xor x960 xor x1511 xor x1607;
a360<=x37 xor x215 xor x809 xor x865 xor x1512 xor x1608;
a361<=x38 xor x216 xor x810 xor x866 xor x1513 xor x1609;
a362<=x39 xor x217 xor x811 xor x867 xor x1514 xor x1610;
a363<=x40 xor x218 xor x812 xor x868 xor x1515 xor x1611;
a364<=x41 xor x219 xor x813 xor x869 xor x1516 xor x1612;
a365<=x42 xor x220 xor x814 xor x870 xor x1517 xor x1613;
a366<=x43 xor x221 xor x815 xor x871 xor x1518 xor x1614;
a367<=x44 xor x222 xor x816 xor x872 xor x1519 xor x1615;
a368<=x45 xor x223 xor x817 xor x873 xor x1520 xor x1616;
a369<=x46 xor x224 xor x818 xor x874 xor x1521 xor x1617;
a370<=x47 xor x225 xor x819 xor x875 xor x1522 xor x1618;
a371<=x48 xor x226 xor x820 xor x876 xor x1523 xor x1619;
a372<=x49 xor x227 xor x821 xor x877 xor x1524 xor x1620;
a373<=x50 xor x228 xor x822 xor x878 xor x1525 xor x1621;
a374<=x51 xor x229 xor x823 xor x879 xor x1526 xor x1622;
a375<=x52 xor x230 xor x824 xor x880 xor x1527 xor x1623;
a376<=x53 xor x231 xor x825 xor x881 xor x1528 xor x1624;
a377<=x54 xor x232 xor x826 xor x882 xor x1529 xor x1625;
a378<=x55 xor x233 xor x827 xor x883 xor x1530 xor x1626;
a379<=x56 xor x234 xor x828 xor x884 xor x1531 xor x1627;
a380<=x57 xor x235 xor x829 xor x885 xor x1532 xor x1628;
a381<=x58 xor x236 xor x830 xor x886 xor x1533 xor x1629;
a382<=x59 xor x237 xor x831 xor x887 xor x1534 xor x1630;
a383<=x60 xor x238 xor x832 xor x888 xor x1535 xor x1631;
a384<=x61 xor x239 xor x833 xor x889 xor x1536 xor x1632;
a385<=x232 xor x661 xor x906 xor x1033 xor x1537 xor x1633;
a386<=x233 xor x662 xor x907 xor x1034 xor x1538 xor x1634;
a387<=x234 xor x663 xor x908 xor x1035 xor x1539 xor x1635;
a388<=x235 xor x664 xor x909 xor x1036 xor x1540 xor x1636;
a389<=x236 xor x665 xor x910 xor x1037 xor x1541 xor x1637;
a390<=x237 xor x666 xor x911 xor x1038 xor x1542 xor x1638;
a391<=x238 xor x667 xor x912 xor x1039 xor x1543 xor x1639;
a392<=x239 xor x668 xor x913 xor x1040 xor x1544 xor x1640;
a393<=x240 xor x669 xor x914 xor x1041 xor x1545 xor x1641;
a394<=x241 xor x670 xor x915 xor x1042 xor x1546 xor x1642;
a395<=x242 xor x671 xor x916 xor x1043 xor x1547 xor x1643;
a396<=x243 xor x672 xor x917 xor x1044 xor x1548 xor x1644;
a397<=x244 xor x577 xor x918 xor x1045 xor x1549 xor x1645;
a398<=x245 xor x578 xor x919 xor x1046 xor x1550 xor x1646;
a399<=x246 xor x579 xor x920 xor x1047 xor x1551 xor x1647;
a400<=x247 xor x580 xor x921 xor x1048 xor x1552 xor x1648;
a401<=x248 xor x581 xor x922 xor x1049 xor x1553 xor x1649;
a402<=x249 xor x582 xor x923 xor x1050 xor x1554 xor x1650;
a403<=x250 xor x583 xor x924 xor x1051 xor x1555 xor x1651;
a404<=x251 xor x584 xor x925 xor x1052 xor x1556 xor x1652;
a405<=x252 xor x585 xor x926 xor x1053 xor x1557 xor x1653;
a406<=x253 xor x586 xor x927 xor x1054 xor x1558 xor x1654;
a407<=x254 xor x587 xor x928 xor x1055 xor x1559 xor x1655;
a408<=x255 xor x588 xor x929 xor x1056 xor x1560 xor x1656;
a409<=x256 xor x589 xor x930 xor x961 xor x1561 xor x1657;
a410<=x257 xor x590 xor x931 xor x962 xor x1562 xor x1658;
a411<=x258 xor x591 xor x932 xor x963 xor x1563 xor x1659;
a412<=x259 xor x592 xor x933 xor x964 xor x1564 xor x1660;
a413<=x260 xor x593 xor x934 xor x965 xor x1565 xor x1661;
a414<=x261 xor x594 xor x935 xor x966 xor x1566 xor x1662;
a415<=x262 xor x595 xor x936 xor x967 xor x1567 xor x1663;
a416<=x263 xor x596 xor x937 xor x968 xor x1568 xor x1664;
a417<=x264 xor x597 xor x938 xor x969 xor x1569 xor x1665;
a418<=x265 xor x598 xor x939 xor x970 xor x1570 xor x1666;
a419<=x266 xor x599 xor x940 xor x971 xor x1571 xor x1667;
a420<=x267 xor x600 xor x941 xor x972 xor x1572 xor x1668;
a421<=x268 xor x601 xor x942 xor x973 xor x1573 xor x1669;
a422<=x269 xor x602 xor x943 xor x974 xor x1574 xor x1670;
a423<=x270 xor x603 xor x944 xor x975 xor x1575 xor x1671;
a424<=x271 xor x604 xor x945 xor x976 xor x1576 xor x1672;
a425<=x272 xor x605 xor x946 xor x977 xor x1577 xor x1673;
a426<=x273 xor x606 xor x947 xor x978 xor x1578 xor x1674;
a427<=x274 xor x607 xor x948 xor x979 xor x1579 xor x1675;
a428<=x275 xor x608 xor x949 xor x980 xor x1580 xor x1676;
a429<=x276 xor x609 xor x950 xor x981 xor x1581 xor x1677;
a430<=x277 xor x610 xor x951 xor x982 xor x1582 xor x1678;
a431<=x278 xor x611 xor x952 xor x983 xor x1583 xor x1679;
a432<=x279 xor x612 xor x953 xor x984 xor x1584 xor x1680;
a433<=x280 xor x613 xor x954 xor x985 xor x1585 xor x1681;
a434<=x281 xor x614 xor x955 xor x986 xor x1586 xor x1682;
a435<=x282 xor x615 xor x956 xor x987 xor x1587 xor x1683;
a436<=x283 xor x616 xor x957 xor x988 xor x1588 xor x1684;
a437<=x284 xor x617 xor x958 xor x989 xor x1589 xor x1685;
a438<=x285 xor x618 xor x959 xor x990 xor x1590 xor x1686;
a439<=x286 xor x619 xor x960 xor x991 xor x1591 xor x1687;
a440<=x287 xor x620 xor x865 xor x992 xor x1592 xor x1688;
a441<=x288 xor x621 xor x866 xor x993 xor x1593 xor x1689;
a442<=x193 xor x622 xor x867 xor x994 xor x1594 xor x1690;
a443<=x194 xor x623 xor x868 xor x995 xor x1595 xor x1691;
a444<=x195 xor x624 xor x869 xor x996 xor x1596 xor x1692;
a445<=x196 xor x625 xor x870 xor x997 xor x1597 xor x1693;
a446<=x197 xor x626 xor x871 xor x998 xor x1598 xor x1694;
a447<=x198 xor x627 xor x872 xor x999 xor x1599 xor x1695;
a448<=x199 xor x628 xor x873 xor x1000 xor x1600 xor x1696;
a449<=x200 xor x629 xor x874 xor x1001 xor x1601 xor x1697;
a450<=x201 xor x630 xor x875 xor x1002 xor x1602 xor x1698;
a451<=x202 xor x631 xor x876 xor x1003 xor x1603 xor x1699;
a452<=x203 xor x632 xor x877 xor x1004 xor x1604 xor x1700;
a453<=x204 xor x633 xor x878 xor x1005 xor x1605 xor x1701;
a454<=x205 xor x634 xor x879 xor x1006 xor x1606 xor x1702;
a455<=x206 xor x635 xor x880 xor x1007 xor x1607 xor x1703;
a456<=x207 xor x636 xor x881 xor x1008 xor x1608 xor x1704;
a457<=x208 xor x637 xor x882 xor x1009 xor x1609 xor x1705;
a458<=x209 xor x638 xor x883 xor x1010 xor x1610 xor x1706;
a459<=x210 xor x639 xor x884 xor x1011 xor x1611 xor x1707;
a460<=x211 xor x640 xor x885 xor x1012 xor x1612 xor x1708;
a461<=x212 xor x641 xor x886 xor x1013 xor x1613 xor x1709;
a462<=x213 xor x642 xor x887 xor x1014 xor x1614 xor x1710;
a463<=x214 xor x643 xor x888 xor x1015 xor x1615 xor x1711;
a464<=x215 xor x644 xor x889 xor x1016 xor x1616 xor x1712;
a465<=x216 xor x645 xor x890 xor x1017 xor x1617 xor x1713;
a466<=x217 xor x646 xor x891 xor x1018 xor x1618 xor x1714;
a467<=x218 xor x647 xor x892 xor x1019 xor x1619 xor x1715;
a468<=x219 xor x648 xor x893 xor x1020 xor x1620 xor x1716;
a469<=x220 xor x649 xor x894 xor x1021 xor x1621 xor x1717;
a470<=x221 xor x650 xor x895 xor x1022 xor x1622 xor x1718;
a471<=x222 xor x651 xor x896 xor x1023 xor x1623 xor x1719;
a472<=x223 xor x652 xor x897 xor x1024 xor x1624 xor x1720;
a473<=x224 xor x653 xor x898 xor x1025 xor x1625 xor x1721;
a474<=x225 xor x654 xor x899 xor x1026 xor x1626 xor x1722;
a475<=x226 xor x655 xor x900 xor x1027 xor x1627 xor x1723;
a476<=x227 xor x656 xor x901 xor x1028 xor x1628 xor x1724;
a477<=x228 xor x657 xor x902 xor x1029 xor x1629 xor x1725;
a478<=x229 xor x658 xor x903 xor x1030 xor x1630 xor x1726;
a479<=x230 xor x659 xor x904 xor x1031 xor x1631 xor x1727;
a480<=x231 xor x660 xor x905 xor x1032 xor x1632 xor x1728;
a481<=x431 xor x521 xor x755 xor x1136 xor x1153 xor x1633 xor x1729;
a482<=x432 xor x522 xor x756 xor x1137 xor x1154 xor x1634 xor x1730;
a483<=x433 xor x523 xor x757 xor x1138 xor x1155 xor x1635 xor x1731;
a484<=x434 xor x524 xor x758 xor x1139 xor x1156 xor x1636 xor x1732;
a485<=x435 xor x525 xor x759 xor x1140 xor x1157 xor x1637 xor x1733;
a486<=x436 xor x526 xor x760 xor x1141 xor x1158 xor x1638 xor x1734;
a487<=x437 xor x527 xor x761 xor x1142 xor x1159 xor x1639 xor x1735;
a488<=x438 xor x528 xor x762 xor x1143 xor x1160 xor x1640 xor x1736;
a489<=x439 xor x529 xor x763 xor x1144 xor x1161 xor x1641 xor x1737;
a490<=x440 xor x530 xor x764 xor x1145 xor x1162 xor x1642 xor x1738;
a491<=x441 xor x531 xor x765 xor x1146 xor x1163 xor x1643 xor x1739;
a492<=x442 xor x532 xor x766 xor x1147 xor x1164 xor x1644 xor x1740;
a493<=x443 xor x533 xor x767 xor x1148 xor x1165 xor x1645 xor x1741;
a494<=x444 xor x534 xor x768 xor x1149 xor x1166 xor x1646 xor x1742;
a495<=x445 xor x535 xor x673 xor x1150 xor x1167 xor x1647 xor x1743;
a496<=x446 xor x536 xor x674 xor x1151 xor x1168 xor x1648 xor x1744;
a497<=x447 xor x537 xor x675 xor x1152 xor x1169 xor x1649 xor x1745;
a498<=x448 xor x538 xor x676 xor x1057 xor x1170 xor x1650 xor x1746;
a499<=x449 xor x539 xor x677 xor x1058 xor x1171 xor x1651 xor x1747;
a500<=x450 xor x540 xor x678 xor x1059 xor x1172 xor x1652 xor x1748;
a501<=x451 xor x541 xor x679 xor x1060 xor x1173 xor x1653 xor x1749;
a502<=x452 xor x542 xor x680 xor x1061 xor x1174 xor x1654 xor x1750;
a503<=x453 xor x543 xor x681 xor x1062 xor x1175 xor x1655 xor x1751;
a504<=x454 xor x544 xor x682 xor x1063 xor x1176 xor x1656 xor x1752;
a505<=x455 xor x545 xor x683 xor x1064 xor x1177 xor x1657 xor x1753;
a506<=x456 xor x546 xor x684 xor x1065 xor x1178 xor x1658 xor x1754;
a507<=x457 xor x547 xor x685 xor x1066 xor x1179 xor x1659 xor x1755;
a508<=x458 xor x548 xor x686 xor x1067 xor x1180 xor x1660 xor x1756;
a509<=x459 xor x549 xor x687 xor x1068 xor x1181 xor x1661 xor x1757;
a510<=x460 xor x550 xor x688 xor x1069 xor x1182 xor x1662 xor x1758;
a511<=x461 xor x551 xor x689 xor x1070 xor x1183 xor x1663 xor x1759;
a512<=x462 xor x552 xor x690 xor x1071 xor x1184 xor x1664 xor x1760;
a513<=x463 xor x553 xor x691 xor x1072 xor x1185 xor x1665 xor x1761;
a514<=x464 xor x554 xor x692 xor x1073 xor x1186 xor x1666 xor x1762;
a515<=x465 xor x555 xor x693 xor x1074 xor x1187 xor x1667 xor x1763;
a516<=x466 xor x556 xor x694 xor x1075 xor x1188 xor x1668 xor x1764;
a517<=x467 xor x557 xor x695 xor x1076 xor x1189 xor x1669 xor x1765;
a518<=x468 xor x558 xor x696 xor x1077 xor x1190 xor x1670 xor x1766;
a519<=x469 xor x559 xor x697 xor x1078 xor x1191 xor x1671 xor x1767;
a520<=x470 xor x560 xor x698 xor x1079 xor x1192 xor x1672 xor x1768;
a521<=x471 xor x561 xor x699 xor x1080 xor x1193 xor x1673 xor x1769;
a522<=x472 xor x562 xor x700 xor x1081 xor x1194 xor x1674 xor x1770;
a523<=x473 xor x563 xor x701 xor x1082 xor x1195 xor x1675 xor x1771;
a524<=x474 xor x564 xor x702 xor x1083 xor x1196 xor x1676 xor x1772;
a525<=x475 xor x565 xor x703 xor x1084 xor x1197 xor x1677 xor x1773;
a526<=x476 xor x566 xor x704 xor x1085 xor x1198 xor x1678 xor x1774;
a527<=x477 xor x567 xor x705 xor x1086 xor x1199 xor x1679 xor x1775;
a528<=x478 xor x568 xor x706 xor x1087 xor x1200 xor x1680 xor x1776;
a529<=x479 xor x569 xor x707 xor x1088 xor x1201 xor x1681 xor x1777;
a530<=x480 xor x570 xor x708 xor x1089 xor x1202 xor x1682 xor x1778;
a531<=x385 xor x571 xor x709 xor x1090 xor x1203 xor x1683 xor x1779;
a532<=x386 xor x572 xor x710 xor x1091 xor x1204 xor x1684 xor x1780;
a533<=x387 xor x573 xor x711 xor x1092 xor x1205 xor x1685 xor x1781;
a534<=x388 xor x574 xor x712 xor x1093 xor x1206 xor x1686 xor x1782;
a535<=x389 xor x575 xor x713 xor x1094 xor x1207 xor x1687 xor x1783;
a536<=x390 xor x576 xor x714 xor x1095 xor x1208 xor x1688 xor x1784;
a537<=x391 xor x481 xor x715 xor x1096 xor x1209 xor x1689 xor x1785;
a538<=x392 xor x482 xor x716 xor x1097 xor x1210 xor x1690 xor x1786;
a539<=x393 xor x483 xor x717 xor x1098 xor x1211 xor x1691 xor x1787;
a540<=x394 xor x484 xor x718 xor x1099 xor x1212 xor x1692 xor x1788;
a541<=x395 xor x485 xor x719 xor x1100 xor x1213 xor x1693 xor x1789;
a542<=x396 xor x486 xor x720 xor x1101 xor x1214 xor x1694 xor x1790;
a543<=x397 xor x487 xor x721 xor x1102 xor x1215 xor x1695 xor x1791;
a544<=x398 xor x488 xor x722 xor x1103 xor x1216 xor x1696 xor x1792;
a545<=x399 xor x489 xor x723 xor x1104 xor x1217 xor x1697 xor x1793;
a546<=x400 xor x490 xor x724 xor x1105 xor x1218 xor x1698 xor x1794;
a547<=x401 xor x491 xor x725 xor x1106 xor x1219 xor x1699 xor x1795;
a548<=x402 xor x492 xor x726 xor x1107 xor x1220 xor x1700 xor x1796;
a549<=x403 xor x493 xor x727 xor x1108 xor x1221 xor x1701 xor x1797;
a550<=x404 xor x494 xor x728 xor x1109 xor x1222 xor x1702 xor x1798;
a551<=x405 xor x495 xor x729 xor x1110 xor x1223 xor x1703 xor x1799;
a552<=x406 xor x496 xor x730 xor x1111 xor x1224 xor x1704 xor x1800;
a553<=x407 xor x497 xor x731 xor x1112 xor x1225 xor x1705 xor x1801;
a554<=x408 xor x498 xor x732 xor x1113 xor x1226 xor x1706 xor x1802;
a555<=x409 xor x499 xor x733 xor x1114 xor x1227 xor x1707 xor x1803;
a556<=x410 xor x500 xor x734 xor x1115 xor x1228 xor x1708 xor x1804;
a557<=x411 xor x501 xor x735 xor x1116 xor x1229 xor x1709 xor x1805;
a558<=x412 xor x502 xor x736 xor x1117 xor x1230 xor x1710 xor x1806;
a559<=x413 xor x503 xor x737 xor x1118 xor x1231 xor x1711 xor x1807;
a560<=x414 xor x504 xor x738 xor x1119 xor x1232 xor x1712 xor x1808;
a561<=x415 xor x505 xor x739 xor x1120 xor x1233 xor x1713 xor x1809;
a562<=x416 xor x506 xor x740 xor x1121 xor x1234 xor x1714 xor x1810;
a563<=x417 xor x507 xor x741 xor x1122 xor x1235 xor x1715 xor x1811;
a564<=x418 xor x508 xor x742 xor x1123 xor x1236 xor x1716 xor x1812;
a565<=x419 xor x509 xor x743 xor x1124 xor x1237 xor x1717 xor x1813;
a566<=x420 xor x510 xor x744 xor x1125 xor x1238 xor x1718 xor x1814;
a567<=x421 xor x511 xor x745 xor x1126 xor x1239 xor x1719 xor x1815;
a568<=x422 xor x512 xor x746 xor x1127 xor x1240 xor x1720 xor x1816;
a569<=x423 xor x513 xor x747 xor x1128 xor x1241 xor x1721 xor x1817;
a570<=x424 xor x514 xor x748 xor x1129 xor x1242 xor x1722 xor x1818;
a571<=x425 xor x515 xor x749 xor x1130 xor x1243 xor x1723 xor x1819;
a572<=x426 xor x516 xor x750 xor x1131 xor x1244 xor x1724 xor x1820;
a573<=x427 xor x517 xor x751 xor x1132 xor x1245 xor x1725 xor x1821;
a574<=x428 xor x518 xor x752 xor x1133 xor x1246 xor x1726 xor x1822;
a575<=x429 xor x519 xor x753 xor x1134 xor x1247 xor x1727 xor x1823;
a576<=x430 xor x520 xor x754 xor x1135 xor x1248 xor x1728 xor x1824;
a577<=x288 xor x342 xor x879 xor x979 xor x1729 xor x1825;
a578<=x193 xor x343 xor x880 xor x980 xor x1730 xor x1826;
a579<=x194 xor x344 xor x881 xor x981 xor x1731 xor x1827;
a580<=x195 xor x345 xor x882 xor x982 xor x1732 xor x1828;
a581<=x196 xor x346 xor x883 xor x983 xor x1733 xor x1829;
a582<=x197 xor x347 xor x884 xor x984 xor x1734 xor x1830;
a583<=x198 xor x348 xor x885 xor x985 xor x1735 xor x1831;
a584<=x199 xor x349 xor x886 xor x986 xor x1736 xor x1832;
a585<=x200 xor x350 xor x887 xor x987 xor x1737 xor x1833;
a586<=x201 xor x351 xor x888 xor x988 xor x1738 xor x1834;
a587<=x202 xor x352 xor x889 xor x989 xor x1739 xor x1835;
a588<=x203 xor x353 xor x890 xor x990 xor x1740 xor x1836;
a589<=x204 xor x354 xor x891 xor x991 xor x1741 xor x1837;
a590<=x205 xor x355 xor x892 xor x992 xor x1742 xor x1838;
a591<=x206 xor x356 xor x893 xor x993 xor x1743 xor x1839;
a592<=x207 xor x357 xor x894 xor x994 xor x1744 xor x1840;
a593<=x208 xor x358 xor x895 xor x995 xor x1745 xor x1841;
a594<=x209 xor x359 xor x896 xor x996 xor x1746 xor x1842;
a595<=x210 xor x360 xor x897 xor x997 xor x1747 xor x1843;
a596<=x211 xor x361 xor x898 xor x998 xor x1748 xor x1844;
a597<=x212 xor x362 xor x899 xor x999 xor x1749 xor x1845;
a598<=x213 xor x363 xor x900 xor x1000 xor x1750 xor x1846;
a599<=x214 xor x364 xor x901 xor x1001 xor x1751 xor x1847;
a600<=x215 xor x365 xor x902 xor x1002 xor x1752 xor x1848;
a601<=x216 xor x366 xor x903 xor x1003 xor x1753 xor x1849;
a602<=x217 xor x367 xor x904 xor x1004 xor x1754 xor x1850;
a603<=x218 xor x368 xor x905 xor x1005 xor x1755 xor x1851;
a604<=x219 xor x369 xor x906 xor x1006 xor x1756 xor x1852;
a605<=x220 xor x370 xor x907 xor x1007 xor x1757 xor x1853;
a606<=x221 xor x371 xor x908 xor x1008 xor x1758 xor x1854;
a607<=x222 xor x372 xor x909 xor x1009 xor x1759 xor x1855;
a608<=x223 xor x373 xor x910 xor x1010 xor x1760 xor x1856;
a609<=x224 xor x374 xor x911 xor x1011 xor x1761 xor x1857;
a610<=x225 xor x375 xor x912 xor x1012 xor x1762 xor x1858;
a611<=x226 xor x376 xor x913 xor x1013 xor x1763 xor x1859;
a612<=x227 xor x377 xor x914 xor x1014 xor x1764 xor x1860;
a613<=x228 xor x378 xor x915 xor x1015 xor x1765 xor x1861;
a614<=x229 xor x379 xor x916 xor x1016 xor x1766 xor x1862;
a615<=x230 xor x380 xor x917 xor x1017 xor x1767 xor x1863;
a616<=x231 xor x381 xor x918 xor x1018 xor x1768 xor x1864;
a617<=x232 xor x382 xor x919 xor x1019 xor x1769 xor x1865;
a618<=x233 xor x383 xor x920 xor x1020 xor x1770 xor x1866;
a619<=x234 xor x384 xor x921 xor x1021 xor x1771 xor x1867;
a620<=x235 xor x289 xor x922 xor x1022 xor x1772 xor x1868;
a621<=x236 xor x290 xor x923 xor x1023 xor x1773 xor x1869;
a622<=x237 xor x291 xor x924 xor x1024 xor x1774 xor x1870;
a623<=x238 xor x292 xor x925 xor x1025 xor x1775 xor x1871;
a624<=x239 xor x293 xor x926 xor x1026 xor x1776 xor x1872;
a625<=x240 xor x294 xor x927 xor x1027 xor x1777 xor x1873;
a626<=x241 xor x295 xor x928 xor x1028 xor x1778 xor x1874;
a627<=x242 xor x296 xor x929 xor x1029 xor x1779 xor x1875;
a628<=x243 xor x297 xor x930 xor x1030 xor x1780 xor x1876;
a629<=x244 xor x298 xor x931 xor x1031 xor x1781 xor x1877;
a630<=x245 xor x299 xor x932 xor x1032 xor x1782 xor x1878;
a631<=x246 xor x300 xor x933 xor x1033 xor x1783 xor x1879;
a632<=x247 xor x301 xor x934 xor x1034 xor x1784 xor x1880;
a633<=x248 xor x302 xor x935 xor x1035 xor x1785 xor x1881;
a634<=x249 xor x303 xor x936 xor x1036 xor x1786 xor x1882;
a635<=x250 xor x304 xor x937 xor x1037 xor x1787 xor x1883;
a636<=x251 xor x305 xor x938 xor x1038 xor x1788 xor x1884;
a637<=x252 xor x306 xor x939 xor x1039 xor x1789 xor x1885;
a638<=x253 xor x307 xor x940 xor x1040 xor x1790 xor x1886;
a639<=x254 xor x308 xor x941 xor x1041 xor x1791 xor x1887;
a640<=x255 xor x309 xor x942 xor x1042 xor x1792 xor x1888;
a641<=x256 xor x310 xor x943 xor x1043 xor x1793 xor x1889;
a642<=x257 xor x311 xor x944 xor x1044 xor x1794 xor x1890;
a643<=x258 xor x312 xor x945 xor x1045 xor x1795 xor x1891;
a644<=x259 xor x313 xor x946 xor x1046 xor x1796 xor x1892;
a645<=x260 xor x314 xor x947 xor x1047 xor x1797 xor x1893;
a646<=x261 xor x315 xor x948 xor x1048 xor x1798 xor x1894;
a647<=x262 xor x316 xor x949 xor x1049 xor x1799 xor x1895;
a648<=x263 xor x317 xor x950 xor x1050 xor x1800 xor x1896;
a649<=x264 xor x318 xor x951 xor x1051 xor x1801 xor x1897;
a650<=x265 xor x319 xor x952 xor x1052 xor x1802 xor x1898;
a651<=x266 xor x320 xor x953 xor x1053 xor x1803 xor x1899;
a652<=x267 xor x321 xor x954 xor x1054 xor x1804 xor x1900;
a653<=x268 xor x322 xor x955 xor x1055 xor x1805 xor x1901;
a654<=x269 xor x323 xor x956 xor x1056 xor x1806 xor x1902;
a655<=x270 xor x324 xor x957 xor x961 xor x1807 xor x1903;
a656<=x271 xor x325 xor x958 xor x962 xor x1808 xor x1904;
a657<=x272 xor x326 xor x959 xor x963 xor x1809 xor x1905;
a658<=x273 xor x327 xor x960 xor x964 xor x1810 xor x1906;
a659<=x274 xor x328 xor x865 xor x965 xor x1811 xor x1907;
a660<=x275 xor x329 xor x866 xor x966 xor x1812 xor x1908;
a661<=x276 xor x330 xor x867 xor x967 xor x1813 xor x1909;
a662<=x277 xor x331 xor x868 xor x968 xor x1814 xor x1910;
a663<=x278 xor x332 xor x869 xor x969 xor x1815 xor x1911;
a664<=x279 xor x333 xor x870 xor x970 xor x1816 xor x1912;
a665<=x280 xor x334 xor x871 xor x971 xor x1817 xor x1913;
a666<=x281 xor x335 xor x872 xor x972 xor x1818 xor x1914;
a667<=x282 xor x336 xor x873 xor x973 xor x1819 xor x1915;
a668<=x283 xor x337 xor x874 xor x974 xor x1820 xor x1916;
a669<=x284 xor x338 xor x875 xor x975 xor x1821 xor x1917;
a670<=x285 xor x339 xor x876 xor x976 xor x1822 xor x1918;
a671<=x286 xor x340 xor x877 xor x977 xor x1823 xor x1919;
a672<=x287 xor x341 xor x878 xor x978 xor x1824 xor x1920;
a673<=x108 xor x266 xor x579 xor x912 xor x1825 xor x1921;
a674<=x109 xor x267 xor x580 xor x913 xor x1826 xor x1922;
a675<=x110 xor x268 xor x581 xor x914 xor x1827 xor x1923;
a676<=x111 xor x269 xor x582 xor x915 xor x1828 xor x1924;
a677<=x112 xor x270 xor x583 xor x916 xor x1829 xor x1925;
a678<=x113 xor x271 xor x584 xor x917 xor x1830 xor x1926;
a679<=x114 xor x272 xor x585 xor x918 xor x1831 xor x1927;
a680<=x115 xor x273 xor x586 xor x919 xor x1832 xor x1928;
a681<=x116 xor x274 xor x587 xor x920 xor x1833 xor x1929;
a682<=x117 xor x275 xor x588 xor x921 xor x1834 xor x1930;
a683<=x118 xor x276 xor x589 xor x922 xor x1835 xor x1931;
a684<=x119 xor x277 xor x590 xor x923 xor x1836 xor x1932;
a685<=x120 xor x278 xor x591 xor x924 xor x1837 xor x1933;
a686<=x121 xor x279 xor x592 xor x925 xor x1838 xor x1934;
a687<=x122 xor x280 xor x593 xor x926 xor x1839 xor x1935;
a688<=x123 xor x281 xor x594 xor x927 xor x1840 xor x1936;
a689<=x124 xor x282 xor x595 xor x928 xor x1841 xor x1937;
a690<=x125 xor x283 xor x596 xor x929 xor x1842 xor x1938;
a691<=x126 xor x284 xor x597 xor x930 xor x1843 xor x1939;
a692<=x127 xor x285 xor x598 xor x931 xor x1844 xor x1940;
a693<=x128 xor x286 xor x599 xor x932 xor x1845 xor x1941;
a694<=x129 xor x287 xor x600 xor x933 xor x1846 xor x1942;
a695<=x130 xor x288 xor x601 xor x934 xor x1847 xor x1943;
a696<=x131 xor x193 xor x602 xor x935 xor x1848 xor x1944;
a697<=x132 xor x194 xor x603 xor x936 xor x1849 xor x1945;
a698<=x133 xor x195 xor x604 xor x937 xor x1850 xor x1946;
a699<=x134 xor x196 xor x605 xor x938 xor x1851 xor x1947;
a700<=x135 xor x197 xor x606 xor x939 xor x1852 xor x1948;
a701<=x136 xor x198 xor x607 xor x940 xor x1853 xor x1949;
a702<=x137 xor x199 xor x608 xor x941 xor x1854 xor x1950;
a703<=x138 xor x200 xor x609 xor x942 xor x1855 xor x1951;
a704<=x139 xor x201 xor x610 xor x943 xor x1856 xor x1952;
a705<=x140 xor x202 xor x611 xor x944 xor x1857 xor x1953;
a706<=x141 xor x203 xor x612 xor x945 xor x1858 xor x1954;
a707<=x142 xor x204 xor x613 xor x946 xor x1859 xor x1955;
a708<=x143 xor x205 xor x614 xor x947 xor x1860 xor x1956;
a709<=x144 xor x206 xor x615 xor x948 xor x1861 xor x1957;
a710<=x145 xor x207 xor x616 xor x949 xor x1862 xor x1958;
a711<=x146 xor x208 xor x617 xor x950 xor x1863 xor x1959;
a712<=x147 xor x209 xor x618 xor x951 xor x1864 xor x1960;
a713<=x148 xor x210 xor x619 xor x952 xor x1865 xor x1961;
a714<=x149 xor x211 xor x620 xor x953 xor x1866 xor x1962;
a715<=x150 xor x212 xor x621 xor x954 xor x1867 xor x1963;
a716<=x151 xor x213 xor x622 xor x955 xor x1868 xor x1964;
a717<=x152 xor x214 xor x623 xor x956 xor x1869 xor x1965;
a718<=x153 xor x215 xor x624 xor x957 xor x1870 xor x1966;
a719<=x154 xor x216 xor x625 xor x958 xor x1871 xor x1967;
a720<=x155 xor x217 xor x626 xor x959 xor x1872 xor x1968;
a721<=x156 xor x218 xor x627 xor x960 xor x1873 xor x1969;
a722<=x157 xor x219 xor x628 xor x865 xor x1874 xor x1970;
a723<=x158 xor x220 xor x629 xor x866 xor x1875 xor x1971;
a724<=x159 xor x221 xor x630 xor x867 xor x1876 xor x1972;
a725<=x160 xor x222 xor x631 xor x868 xor x1877 xor x1973;
a726<=x161 xor x223 xor x632 xor x869 xor x1878 xor x1974;
a727<=x162 xor x224 xor x633 xor x870 xor x1879 xor x1975;
a728<=x163 xor x225 xor x634 xor x871 xor x1880 xor x1976;
a729<=x164 xor x226 xor x635 xor x872 xor x1881 xor x1977;
a730<=x165 xor x227 xor x636 xor x873 xor x1882 xor x1978;
a731<=x166 xor x228 xor x637 xor x874 xor x1883 xor x1979;
a732<=x167 xor x229 xor x638 xor x875 xor x1884 xor x1980;
a733<=x168 xor x230 xor x639 xor x876 xor x1885 xor x1981;
a734<=x169 xor x231 xor x640 xor x877 xor x1886 xor x1982;
a735<=x170 xor x232 xor x641 xor x878 xor x1887 xor x1983;
a736<=x171 xor x233 xor x642 xor x879 xor x1888 xor x1984;
a737<=x172 xor x234 xor x643 xor x880 xor x1889 xor x1985;
a738<=x173 xor x235 xor x644 xor x881 xor x1890 xor x1986;
a739<=x174 xor x236 xor x645 xor x882 xor x1891 xor x1987;
a740<=x175 xor x237 xor x646 xor x883 xor x1892 xor x1988;
a741<=x176 xor x238 xor x647 xor x884 xor x1893 xor x1989;
a742<=x177 xor x239 xor x648 xor x885 xor x1894 xor x1990;
a743<=x178 xor x240 xor x649 xor x886 xor x1895 xor x1991;
a744<=x179 xor x241 xor x650 xor x887 xor x1896 xor x1992;
a745<=x180 xor x242 xor x651 xor x888 xor x1897 xor x1993;
a746<=x181 xor x243 xor x652 xor x889 xor x1898 xor x1994;
a747<=x182 xor x244 xor x653 xor x890 xor x1899 xor x1995;
a748<=x183 xor x245 xor x654 xor x891 xor x1900 xor x1996;
a749<=x184 xor x246 xor x655 xor x892 xor x1901 xor x1997;
a750<=x185 xor x247 xor x656 xor x893 xor x1902 xor x1998;
a751<=x186 xor x248 xor x657 xor x894 xor x1903 xor x1999;
a752<=x187 xor x249 xor x658 xor x895 xor x1904 xor x2000;
a753<=x188 xor x250 xor x659 xor x896 xor x1905 xor x2001;
a754<=x189 xor x251 xor x660 xor x897 xor x1906 xor x2002;
a755<=x190 xor x252 xor x661 xor x898 xor x1907 xor x2003;
a756<=x191 xor x253 xor x662 xor x899 xor x1908 xor x2004;
a757<=x192 xor x254 xor x663 xor x900 xor x1909 xor x2005;
a758<=x97 xor x255 xor x664 xor x901 xor x1910 xor x2006;
a759<=x98 xor x256 xor x665 xor x902 xor x1911 xor x2007;
a760<=x99 xor x257 xor x666 xor x903 xor x1912 xor x2008;
a761<=x100 xor x258 xor x667 xor x904 xor x1913 xor x2009;
a762<=x101 xor x259 xor x668 xor x905 xor x1914 xor x2010;
a763<=x102 xor x260 xor x669 xor x906 xor x1915 xor x2011;
a764<=x103 xor x261 xor x670 xor x907 xor x1916 xor x2012;
a765<=x104 xor x262 xor x671 xor x908 xor x1917 xor x2013;
a766<=x105 xor x263 xor x672 xor x909 xor x1918 xor x2014;
a767<=x106 xor x264 xor x577 xor x910 xor x1919 xor x2015;
a768<=x107 xor x265 xor x578 xor x911 xor x1920 xor x2016;
a769<=x13 xor x468 xor x505 xor x716 xor x1108 xor x1921 xor x2017;
a770<=x14 xor x469 xor x506 xor x717 xor x1109 xor x1922 xor x2018;
a771<=x15 xor x470 xor x507 xor x718 xor x1110 xor x1923 xor x2019;
a772<=x16 xor x471 xor x508 xor x719 xor x1111 xor x1924 xor x2020;
a773<=x17 xor x472 xor x509 xor x720 xor x1112 xor x1925 xor x2021;
a774<=x18 xor x473 xor x510 xor x721 xor x1113 xor x1926 xor x2022;
a775<=x19 xor x474 xor x511 xor x722 xor x1114 xor x1927 xor x2023;
a776<=x20 xor x475 xor x512 xor x723 xor x1115 xor x1928 xor x2024;
a777<=x21 xor x476 xor x513 xor x724 xor x1116 xor x1929 xor x2025;
a778<=x22 xor x477 xor x514 xor x725 xor x1117 xor x1930 xor x2026;
a779<=x23 xor x478 xor x515 xor x726 xor x1118 xor x1931 xor x2027;
a780<=x24 xor x479 xor x516 xor x727 xor x1119 xor x1932 xor x2028;
a781<=x25 xor x480 xor x517 xor x728 xor x1120 xor x1933 xor x2029;
a782<=x26 xor x385 xor x518 xor x729 xor x1121 xor x1934 xor x2030;
a783<=x27 xor x386 xor x519 xor x730 xor x1122 xor x1935 xor x2031;
a784<=x28 xor x387 xor x520 xor x731 xor x1123 xor x1936 xor x2032;
a785<=x29 xor x388 xor x521 xor x732 xor x1124 xor x1937 xor x2033;
a786<=x30 xor x389 xor x522 xor x733 xor x1125 xor x1938 xor x2034;
a787<=x31 xor x390 xor x523 xor x734 xor x1126 xor x1939 xor x2035;
a788<=x32 xor x391 xor x524 xor x735 xor x1127 xor x1940 xor x2036;
a789<=x33 xor x392 xor x525 xor x736 xor x1128 xor x1941 xor x2037;
a790<=x34 xor x393 xor x526 xor x737 xor x1129 xor x1942 xor x2038;
a791<=x35 xor x394 xor x527 xor x738 xor x1130 xor x1943 xor x2039;
a792<=x36 xor x395 xor x528 xor x739 xor x1131 xor x1944 xor x2040;
a793<=x37 xor x396 xor x529 xor x740 xor x1132 xor x1945 xor x2041;
a794<=x38 xor x397 xor x530 xor x741 xor x1133 xor x1946 xor x2042;
a795<=x39 xor x398 xor x531 xor x742 xor x1134 xor x1947 xor x2043;
a796<=x40 xor x399 xor x532 xor x743 xor x1135 xor x1948 xor x2044;
a797<=x41 xor x400 xor x533 xor x744 xor x1136 xor x1949 xor x2045;
a798<=x42 xor x401 xor x534 xor x745 xor x1137 xor x1950 xor x2046;
a799<=x43 xor x402 xor x535 xor x746 xor x1138 xor x1951 xor x2047;
a800<=x44 xor x403 xor x536 xor x747 xor x1139 xor x1952 xor x2048;
a801<=x45 xor x404 xor x537 xor x748 xor x1140 xor x1953 xor x2049;
a802<=x46 xor x405 xor x538 xor x749 xor x1141 xor x1954 xor x2050;
a803<=x47 xor x406 xor x539 xor x750 xor x1142 xor x1955 xor x2051;
a804<=x48 xor x407 xor x540 xor x751 xor x1143 xor x1956 xor x2052;
a805<=x49 xor x408 xor x541 xor x752 xor x1144 xor x1957 xor x2053;
a806<=x50 xor x409 xor x542 xor x753 xor x1145 xor x1958 xor x2054;
a807<=x51 xor x410 xor x543 xor x754 xor x1146 xor x1959 xor x2055;
a808<=x52 xor x411 xor x544 xor x755 xor x1147 xor x1960 xor x2056;
a809<=x53 xor x412 xor x545 xor x756 xor x1148 xor x1961 xor x2057;
a810<=x54 xor x413 xor x546 xor x757 xor x1149 xor x1962 xor x2058;
a811<=x55 xor x414 xor x547 xor x758 xor x1150 xor x1963 xor x2059;
a812<=x56 xor x415 xor x548 xor x759 xor x1151 xor x1964 xor x2060;
a813<=x57 xor x416 xor x549 xor x760 xor x1152 xor x1965 xor x2061;
a814<=x58 xor x417 xor x550 xor x761 xor x1057 xor x1966 xor x2062;
a815<=x59 xor x418 xor x551 xor x762 xor x1058 xor x1967 xor x2063;
a816<=x60 xor x419 xor x552 xor x763 xor x1059 xor x1968 xor x2064;
a817<=x61 xor x420 xor x553 xor x764 xor x1060 xor x1969 xor x2065;
a818<=x62 xor x421 xor x554 xor x765 xor x1061 xor x1970 xor x2066;
a819<=x63 xor x422 xor x555 xor x766 xor x1062 xor x1971 xor x2067;
a820<=x64 xor x423 xor x556 xor x767 xor x1063 xor x1972 xor x2068;
a821<=x65 xor x424 xor x557 xor x768 xor x1064 xor x1973 xor x2069;
a822<=x66 xor x425 xor x558 xor x673 xor x1065 xor x1974 xor x2070;
a823<=x67 xor x426 xor x559 xor x674 xor x1066 xor x1975 xor x2071;
a824<=x68 xor x427 xor x560 xor x675 xor x1067 xor x1976 xor x2072;
a825<=x69 xor x428 xor x561 xor x676 xor x1068 xor x1977 xor x2073;
a826<=x70 xor x429 xor x562 xor x677 xor x1069 xor x1978 xor x2074;
a827<=x71 xor x430 xor x563 xor x678 xor x1070 xor x1979 xor x2075;
a828<=x72 xor x431 xor x564 xor x679 xor x1071 xor x1980 xor x2076;
a829<=x73 xor x432 xor x565 xor x680 xor x1072 xor x1981 xor x2077;
a830<=x74 xor x433 xor x566 xor x681 xor x1073 xor x1982 xor x2078;
a831<=x75 xor x434 xor x567 xor x682 xor x1074 xor x1983 xor x2079;
a832<=x76 xor x435 xor x568 xor x683 xor x1075 xor x1984 xor x2080;
a833<=x77 xor x436 xor x569 xor x684 xor x1076 xor x1985 xor x2081;
a834<=x78 xor x437 xor x570 xor x685 xor x1077 xor x1986 xor x2082;
a835<=x79 xor x438 xor x571 xor x686 xor x1078 xor x1987 xor x2083;
a836<=x80 xor x439 xor x572 xor x687 xor x1079 xor x1988 xor x2084;
a837<=x81 xor x440 xor x573 xor x688 xor x1080 xor x1989 xor x2085;
a838<=x82 xor x441 xor x574 xor x689 xor x1081 xor x1990 xor x2086;
a839<=x83 xor x442 xor x575 xor x690 xor x1082 xor x1991 xor x2087;
a840<=x84 xor x443 xor x576 xor x691 xor x1083 xor x1992 xor x2088;
a841<=x85 xor x444 xor x481 xor x692 xor x1084 xor x1993 xor x2089;
a842<=x86 xor x445 xor x482 xor x693 xor x1085 xor x1994 xor x2090;
a843<=x87 xor x446 xor x483 xor x694 xor x1086 xor x1995 xor x2091;
a844<=x88 xor x447 xor x484 xor x695 xor x1087 xor x1996 xor x2092;
a845<=x89 xor x448 xor x485 xor x696 xor x1088 xor x1997 xor x2093;
a846<=x90 xor x449 xor x486 xor x697 xor x1089 xor x1998 xor x2094;
a847<=x91 xor x450 xor x487 xor x698 xor x1090 xor x1999 xor x2095;
a848<=x92 xor x451 xor x488 xor x699 xor x1091 xor x2000 xor x2096;
a849<=x93 xor x452 xor x489 xor x700 xor x1092 xor x2001 xor x2097;
a850<=x94 xor x453 xor x490 xor x701 xor x1093 xor x2002 xor x2098;
a851<=x95 xor x454 xor x491 xor x702 xor x1094 xor x2003 xor x2099;
a852<=x96 xor x455 xor x492 xor x703 xor x1095 xor x2004 xor x2100;
a853<=x1 xor x456 xor x493 xor x704 xor x1096 xor x2005 xor x2101;
a854<=x2 xor x457 xor x494 xor x705 xor x1097 xor x2006 xor x2102;
a855<=x3 xor x458 xor x495 xor x706 xor x1098 xor x2007 xor x2103;
a856<=x4 xor x459 xor x496 xor x707 xor x1099 xor x2008 xor x2104;
a857<=x5 xor x460 xor x497 xor x708 xor x1100 xor x2009 xor x2105;
a858<=x6 xor x461 xor x498 xor x709 xor x1101 xor x2010 xor x2106;
a859<=x7 xor x462 xor x499 xor x710 xor x1102 xor x2011 xor x2107;
a860<=x8 xor x463 xor x500 xor x711 xor x1103 xor x2012 xor x2108;
a861<=x9 xor x464 xor x501 xor x712 xor x1104 xor x2013 xor x2109;
a862<=x10 xor x465 xor x502 xor x713 xor x1105 xor x2014 xor x2110;
a863<=x11 xor x466 xor x503 xor x714 xor x1106 xor x2015 xor x2111;
a864<=x12 xor x467 xor x504 xor x715 xor x1107 xor x2016 xor x2112;
a865<=x575 xor x732 xor x1031 xor x1129 xor x2017 xor x2113;
a866<=x576 xor x733 xor x1032 xor x1130 xor x2018 xor x2114;
a867<=x481 xor x734 xor x1033 xor x1131 xor x2019 xor x2115;
a868<=x482 xor x735 xor x1034 xor x1132 xor x2020 xor x2116;
a869<=x483 xor x736 xor x1035 xor x1133 xor x2021 xor x2117;
a870<=x484 xor x737 xor x1036 xor x1134 xor x2022 xor x2118;
a871<=x485 xor x738 xor x1037 xor x1135 xor x2023 xor x2119;
a872<=x486 xor x739 xor x1038 xor x1136 xor x2024 xor x2120;
a873<=x487 xor x740 xor x1039 xor x1137 xor x2025 xor x2121;
a874<=x488 xor x741 xor x1040 xor x1138 xor x2026 xor x2122;
a875<=x489 xor x742 xor x1041 xor x1139 xor x2027 xor x2123;
a876<=x490 xor x743 xor x1042 xor x1140 xor x2028 xor x2124;
a877<=x491 xor x744 xor x1043 xor x1141 xor x2029 xor x2125;
a878<=x492 xor x745 xor x1044 xor x1142 xor x2030 xor x2126;
a879<=x493 xor x746 xor x1045 xor x1143 xor x2031 xor x2127;
a880<=x494 xor x747 xor x1046 xor x1144 xor x2032 xor x2128;
a881<=x495 xor x748 xor x1047 xor x1145 xor x2033 xor x2129;
a882<=x496 xor x749 xor x1048 xor x1146 xor x2034 xor x2130;
a883<=x497 xor x750 xor x1049 xor x1147 xor x2035 xor x2131;
a884<=x498 xor x751 xor x1050 xor x1148 xor x2036 xor x2132;
a885<=x499 xor x752 xor x1051 xor x1149 xor x2037 xor x2133;
a886<=x500 xor x753 xor x1052 xor x1150 xor x2038 xor x2134;
a887<=x501 xor x754 xor x1053 xor x1151 xor x2039 xor x2135;
a888<=x502 xor x755 xor x1054 xor x1152 xor x2040 xor x2136;
a889<=x503 xor x756 xor x1055 xor x1057 xor x2041 xor x2137;
a890<=x504 xor x757 xor x1056 xor x1058 xor x2042 xor x2138;
a891<=x505 xor x758 xor x961 xor x1059 xor x2043 xor x2139;
a892<=x506 xor x759 xor x962 xor x1060 xor x2044 xor x2140;
a893<=x507 xor x760 xor x963 xor x1061 xor x2045 xor x2141;
a894<=x508 xor x761 xor x964 xor x1062 xor x2046 xor x2142;
a895<=x509 xor x762 xor x965 xor x1063 xor x2047 xor x2143;
a896<=x510 xor x763 xor x966 xor x1064 xor x2048 xor x2144;
a897<=x511 xor x764 xor x967 xor x1065 xor x2049 xor x2145;
a898<=x512 xor x765 xor x968 xor x1066 xor x2050 xor x2146;
a899<=x513 xor x766 xor x969 xor x1067 xor x2051 xor x2147;
a900<=x514 xor x767 xor x970 xor x1068 xor x2052 xor x2148;
a901<=x515 xor x768 xor x971 xor x1069 xor x2053 xor x2149;
a902<=x516 xor x673 xor x972 xor x1070 xor x2054 xor x2150;
a903<=x517 xor x674 xor x973 xor x1071 xor x2055 xor x2151;
a904<=x518 xor x675 xor x974 xor x1072 xor x2056 xor x2152;
a905<=x519 xor x676 xor x975 xor x1073 xor x2057 xor x2153;
a906<=x520 xor x677 xor x976 xor x1074 xor x2058 xor x2154;
a907<=x521 xor x678 xor x977 xor x1075 xor x2059 xor x2155;
a908<=x522 xor x679 xor x978 xor x1076 xor x2060 xor x2156;
a909<=x523 xor x680 xor x979 xor x1077 xor x2061 xor x2157;
a910<=x524 xor x681 xor x980 xor x1078 xor x2062 xor x2158;
a911<=x525 xor x682 xor x981 xor x1079 xor x2063 xor x2159;
a912<=x526 xor x683 xor x982 xor x1080 xor x2064 xor x2160;
a913<=x527 xor x684 xor x983 xor x1081 xor x2065 xor x2161;
a914<=x528 xor x685 xor x984 xor x1082 xor x2066 xor x2162;
a915<=x529 xor x686 xor x985 xor x1083 xor x2067 xor x2163;
a916<=x530 xor x687 xor x986 xor x1084 xor x2068 xor x2164;
a917<=x531 xor x688 xor x987 xor x1085 xor x2069 xor x2165;
a918<=x532 xor x689 xor x988 xor x1086 xor x2070 xor x2166;
a919<=x533 xor x690 xor x989 xor x1087 xor x2071 xor x2167;
a920<=x534 xor x691 xor x990 xor x1088 xor x2072 xor x2168;
a921<=x535 xor x692 xor x991 xor x1089 xor x2073 xor x2169;
a922<=x536 xor x693 xor x992 xor x1090 xor x2074 xor x2170;
a923<=x537 xor x694 xor x993 xor x1091 xor x2075 xor x2171;
a924<=x538 xor x695 xor x994 xor x1092 xor x2076 xor x2172;
a925<=x539 xor x696 xor x995 xor x1093 xor x2077 xor x2173;
a926<=x540 xor x697 xor x996 xor x1094 xor x2078 xor x2174;
a927<=x541 xor x698 xor x997 xor x1095 xor x2079 xor x2175;
a928<=x542 xor x699 xor x998 xor x1096 xor x2080 xor x2176;
a929<=x543 xor x700 xor x999 xor x1097 xor x2081 xor x2177;
a930<=x544 xor x701 xor x1000 xor x1098 xor x2082 xor x2178;
a931<=x545 xor x702 xor x1001 xor x1099 xor x2083 xor x2179;
a932<=x546 xor x703 xor x1002 xor x1100 xor x2084 xor x2180;
a933<=x547 xor x704 xor x1003 xor x1101 xor x2085 xor x2181;
a934<=x548 xor x705 xor x1004 xor x1102 xor x2086 xor x2182;
a935<=x549 xor x706 xor x1005 xor x1103 xor x2087 xor x2183;
a936<=x550 xor x707 xor x1006 xor x1104 xor x2088 xor x2184;
a937<=x551 xor x708 xor x1007 xor x1105 xor x2089 xor x2185;
a938<=x552 xor x709 xor x1008 xor x1106 xor x2090 xor x2186;
a939<=x553 xor x710 xor x1009 xor x1107 xor x2091 xor x2187;
a940<=x554 xor x711 xor x1010 xor x1108 xor x2092 xor x2188;
a941<=x555 xor x712 xor x1011 xor x1109 xor x2093 xor x2189;
a942<=x556 xor x713 xor x1012 xor x1110 xor x2094 xor x2190;
a943<=x557 xor x714 xor x1013 xor x1111 xor x2095 xor x2191;
a944<=x558 xor x715 xor x1014 xor x1112 xor x2096 xor x2192;
a945<=x559 xor x716 xor x1015 xor x1113 xor x2097 xor x2193;
a946<=x560 xor x717 xor x1016 xor x1114 xor x2098 xor x2194;
a947<=x561 xor x718 xor x1017 xor x1115 xor x2099 xor x2195;
a948<=x562 xor x719 xor x1018 xor x1116 xor x2100 xor x2196;
a949<=x563 xor x720 xor x1019 xor x1117 xor x2101 xor x2197;
a950<=x564 xor x721 xor x1020 xor x1118 xor x2102 xor x2198;
a951<=x565 xor x722 xor x1021 xor x1119 xor x2103 xor x2199;
a952<=x566 xor x723 xor x1022 xor x1120 xor x2104 xor x2200;
a953<=x567 xor x724 xor x1023 xor x1121 xor x2105 xor x2201;
a954<=x568 xor x725 xor x1024 xor x1122 xor x2106 xor x2202;
a955<=x569 xor x726 xor x1025 xor x1123 xor x2107 xor x2203;
a956<=x570 xor x727 xor x1026 xor x1124 xor x2108 xor x2204;
a957<=x571 xor x728 xor x1027 xor x1125 xor x2109 xor x2205;
a958<=x572 xor x729 xor x1028 xor x1126 xor x2110 xor x2206;
a959<=x573 xor x730 xor x1029 xor x1127 xor x2111 xor x2207;
a960<=x574 xor x731 xor x1030 xor x1128 xor x2112 xor x2208;
a961<=x200 xor x354 xor x808 xor x914 xor x2113 xor x2209;
a962<=x201 xor x355 xor x809 xor x915 xor x2114 xor x2210;
a963<=x202 xor x356 xor x810 xor x916 xor x2115 xor x2211;
a964<=x203 xor x357 xor x811 xor x917 xor x2116 xor x2212;
a965<=x204 xor x358 xor x812 xor x918 xor x2117 xor x2213;
a966<=x205 xor x359 xor x813 xor x919 xor x2118 xor x2214;
a967<=x206 xor x360 xor x814 xor x920 xor x2119 xor x2215;
a968<=x207 xor x361 xor x815 xor x921 xor x2120 xor x2216;
a969<=x208 xor x362 xor x816 xor x922 xor x2121 xor x2217;
a970<=x209 xor x363 xor x817 xor x923 xor x2122 xor x2218;
a971<=x210 xor x364 xor x818 xor x924 xor x2123 xor x2219;
a972<=x211 xor x365 xor x819 xor x925 xor x2124 xor x2220;
a973<=x212 xor x366 xor x820 xor x926 xor x2125 xor x2221;
a974<=x213 xor x367 xor x821 xor x927 xor x2126 xor x2222;
a975<=x214 xor x368 xor x822 xor x928 xor x2127 xor x2223;
a976<=x215 xor x369 xor x823 xor x929 xor x2128 xor x2224;
a977<=x216 xor x370 xor x824 xor x930 xor x2129 xor x2225;
a978<=x217 xor x371 xor x825 xor x931 xor x2130 xor x2226;
a979<=x218 xor x372 xor x826 xor x932 xor x2131 xor x2227;
a980<=x219 xor x373 xor x827 xor x933 xor x2132 xor x2228;
a981<=x220 xor x374 xor x828 xor x934 xor x2133 xor x2229;
a982<=x221 xor x375 xor x829 xor x935 xor x2134 xor x2230;
a983<=x222 xor x376 xor x830 xor x936 xor x2135 xor x2231;
a984<=x223 xor x377 xor x831 xor x937 xor x2136 xor x2232;
a985<=x224 xor x378 xor x832 xor x938 xor x2137 xor x2233;
a986<=x225 xor x379 xor x833 xor x939 xor x2138 xor x2234;
a987<=x226 xor x380 xor x834 xor x940 xor x2139 xor x2235;
a988<=x227 xor x381 xor x835 xor x941 xor x2140 xor x2236;
a989<=x228 xor x382 xor x836 xor x942 xor x2141 xor x2237;
a990<=x229 xor x383 xor x837 xor x943 xor x2142 xor x2238;
a991<=x230 xor x384 xor x838 xor x944 xor x2143 xor x2239;
a992<=x231 xor x289 xor x839 xor x945 xor x2144 xor x2240;
a993<=x232 xor x290 xor x840 xor x946 xor x2145 xor x2241;
a994<=x233 xor x291 xor x841 xor x947 xor x2146 xor x2242;
a995<=x234 xor x292 xor x842 xor x948 xor x2147 xor x2243;
a996<=x235 xor x293 xor x843 xor x949 xor x2148 xor x2244;
a997<=x236 xor x294 xor x844 xor x950 xor x2149 xor x2245;
a998<=x237 xor x295 xor x845 xor x951 xor x2150 xor x2246;
a999<=x238 xor x296 xor x846 xor x952 xor x2151 xor x2247;
a1000<=x239 xor x297 xor x847 xor x953 xor x2152 xor x2248;
a1001<=x240 xor x298 xor x848 xor x954 xor x2153 xor x2249;
a1002<=x241 xor x299 xor x849 xor x955 xor x2154 xor x2250;
a1003<=x242 xor x300 xor x850 xor x956 xor x2155 xor x2251;
a1004<=x243 xor x301 xor x851 xor x957 xor x2156 xor x2252;
a1005<=x244 xor x302 xor x852 xor x958 xor x2157 xor x2253;
a1006<=x245 xor x303 xor x853 xor x959 xor x2158 xor x2254;
a1007<=x246 xor x304 xor x854 xor x960 xor x2159 xor x2255;
a1008<=x247 xor x305 xor x855 xor x865 xor x2160 xor x2256;
a1009<=x248 xor x306 xor x856 xor x866 xor x2161 xor x2257;
a1010<=x249 xor x307 xor x857 xor x867 xor x2162 xor x2258;
a1011<=x250 xor x308 xor x858 xor x868 xor x2163 xor x2259;
a1012<=x251 xor x309 xor x859 xor x869 xor x2164 xor x2260;
a1013<=x252 xor x310 xor x860 xor x870 xor x2165 xor x2261;
a1014<=x253 xor x311 xor x861 xor x871 xor x2166 xor x2262;
a1015<=x254 xor x312 xor x862 xor x872 xor x2167 xor x2263;
a1016<=x255 xor x313 xor x863 xor x873 xor x2168 xor x2264;
a1017<=x256 xor x314 xor x864 xor x874 xor x2169 xor x2265;
a1018<=x257 xor x315 xor x769 xor x875 xor x2170 xor x2266;
a1019<=x258 xor x316 xor x770 xor x876 xor x2171 xor x2267;
a1020<=x259 xor x317 xor x771 xor x877 xor x2172 xor x2268;
a1021<=x260 xor x318 xor x772 xor x878 xor x2173 xor x2269;
a1022<=x261 xor x319 xor x773 xor x879 xor x2174 xor x2270;
a1023<=x262 xor x320 xor x774 xor x880 xor x2175 xor x2271;
a1024<=x263 xor x321 xor x775 xor x881 xor x2176 xor x2272;
a1025<=x264 xor x322 xor x776 xor x882 xor x2177 xor x2273;
a1026<=x265 xor x323 xor x777 xor x883 xor x2178 xor x2274;
a1027<=x266 xor x324 xor x778 xor x884 xor x2179 xor x2275;
a1028<=x267 xor x325 xor x779 xor x885 xor x2180 xor x2276;
a1029<=x268 xor x326 xor x780 xor x886 xor x2181 xor x2277;
a1030<=x269 xor x327 xor x781 xor x887 xor x2182 xor x2278;
a1031<=x270 xor x328 xor x782 xor x888 xor x2183 xor x2279;
a1032<=x271 xor x329 xor x783 xor x889 xor x2184 xor x2280;
a1033<=x272 xor x330 xor x784 xor x890 xor x2185 xor x2281;
a1034<=x273 xor x331 xor x785 xor x891 xor x2186 xor x2282;
a1035<=x274 xor x332 xor x786 xor x892 xor x2187 xor x2283;
a1036<=x275 xor x333 xor x787 xor x893 xor x2188 xor x2284;
a1037<=x276 xor x334 xor x788 xor x894 xor x2189 xor x2285;
a1038<=x277 xor x335 xor x789 xor x895 xor x2190 xor x2286;
a1039<=x278 xor x336 xor x790 xor x896 xor x2191 xor x2287;
a1040<=x279 xor x337 xor x791 xor x897 xor x2192 xor x2288;
a1041<=x280 xor x338 xor x792 xor x898 xor x2193 xor x2289;
a1042<=x281 xor x339 xor x793 xor x899 xor x2194 xor x2290;
a1043<=x282 xor x340 xor x794 xor x900 xor x2195 xor x2291;
a1044<=x283 xor x341 xor x795 xor x901 xor x2196 xor x2292;
a1045<=x284 xor x342 xor x796 xor x902 xor x2197 xor x2293;
a1046<=x285 xor x343 xor x797 xor x903 xor x2198 xor x2294;
a1047<=x286 xor x344 xor x798 xor x904 xor x2199 xor x2295;
a1048<=x287 xor x345 xor x799 xor x905 xor x2200 xor x2296;
a1049<=x288 xor x346 xor x800 xor x906 xor x2201 xor x2297;
a1050<=x193 xor x347 xor x801 xor x907 xor x2202 xor x2298;
a1051<=x194 xor x348 xor x802 xor x908 xor x2203 xor x2299;
a1052<=x195 xor x349 xor x803 xor x909 xor x2204 xor x2300;
a1053<=x196 xor x350 xor x804 xor x910 xor x2205 xor x2301;
a1054<=x197 xor x351 xor x805 xor x911 xor x2206 xor x2302;
a1055<=x198 xor x352 xor x806 xor x912 xor x2207 xor x2303;
a1056<=x199 xor x353 xor x807 xor x913 xor x2208 xor x2304;
a1057<=x44 xor x547 xor x714 xor x1083 xor x1160 xor x2209;
a1058<=x45 xor x548 xor x715 xor x1084 xor x1161 xor x2210;
a1059<=x46 xor x549 xor x716 xor x1085 xor x1162 xor x2211;
a1060<=x47 xor x550 xor x717 xor x1086 xor x1163 xor x2212;
a1061<=x48 xor x551 xor x718 xor x1087 xor x1164 xor x2213;
a1062<=x49 xor x552 xor x719 xor x1088 xor x1165 xor x2214;
a1063<=x50 xor x553 xor x720 xor x1089 xor x1166 xor x2215;
a1064<=x51 xor x554 xor x721 xor x1090 xor x1167 xor x2216;
a1065<=x52 xor x555 xor x722 xor x1091 xor x1168 xor x2217;
a1066<=x53 xor x556 xor x723 xor x1092 xor x1169 xor x2218;
a1067<=x54 xor x557 xor x724 xor x1093 xor x1170 xor x2219;
a1068<=x55 xor x558 xor x725 xor x1094 xor x1171 xor x2220;
a1069<=x56 xor x559 xor x726 xor x1095 xor x1172 xor x2221;
a1070<=x57 xor x560 xor x727 xor x1096 xor x1173 xor x2222;
a1071<=x58 xor x561 xor x728 xor x1097 xor x1174 xor x2223;
a1072<=x59 xor x562 xor x729 xor x1098 xor x1175 xor x2224;
a1073<=x60 xor x563 xor x730 xor x1099 xor x1176 xor x2225;
a1074<=x61 xor x564 xor x731 xor x1100 xor x1177 xor x2226;
a1075<=x62 xor x565 xor x732 xor x1101 xor x1178 xor x2227;
a1076<=x63 xor x566 xor x733 xor x1102 xor x1179 xor x2228;
a1077<=x64 xor x567 xor x734 xor x1103 xor x1180 xor x2229;
a1078<=x65 xor x568 xor x735 xor x1104 xor x1181 xor x2230;
a1079<=x66 xor x569 xor x736 xor x1105 xor x1182 xor x2231;
a1080<=x67 xor x570 xor x737 xor x1106 xor x1183 xor x2232;
a1081<=x68 xor x571 xor x738 xor x1107 xor x1184 xor x2233;
a1082<=x69 xor x572 xor x739 xor x1108 xor x1185 xor x2234;
a1083<=x70 xor x573 xor x740 xor x1109 xor x1186 xor x2235;
a1084<=x71 xor x574 xor x741 xor x1110 xor x1187 xor x2236;
a1085<=x72 xor x575 xor x742 xor x1111 xor x1188 xor x2237;
a1086<=x73 xor x576 xor x743 xor x1112 xor x1189 xor x2238;
a1087<=x74 xor x481 xor x744 xor x1113 xor x1190 xor x2239;
a1088<=x75 xor x482 xor x745 xor x1114 xor x1191 xor x2240;
a1089<=x76 xor x483 xor x746 xor x1115 xor x1192 xor x2241;
a1090<=x77 xor x484 xor x747 xor x1116 xor x1193 xor x2242;
a1091<=x78 xor x485 xor x748 xor x1117 xor x1194 xor x2243;
a1092<=x79 xor x486 xor x749 xor x1118 xor x1195 xor x2244;
a1093<=x80 xor x487 xor x750 xor x1119 xor x1196 xor x2245;
a1094<=x81 xor x488 xor x751 xor x1120 xor x1197 xor x2246;
a1095<=x82 xor x489 xor x752 xor x1121 xor x1198 xor x2247;
a1096<=x83 xor x490 xor x753 xor x1122 xor x1199 xor x2248;
a1097<=x84 xor x491 xor x754 xor x1123 xor x1200 xor x2249;
a1098<=x85 xor x492 xor x755 xor x1124 xor x1201 xor x2250;
a1099<=x86 xor x493 xor x756 xor x1125 xor x1202 xor x2251;
a1100<=x87 xor x494 xor x757 xor x1126 xor x1203 xor x2252;
a1101<=x88 xor x495 xor x758 xor x1127 xor x1204 xor x2253;
a1102<=x89 xor x496 xor x759 xor x1128 xor x1205 xor x2254;
a1103<=x90 xor x497 xor x760 xor x1129 xor x1206 xor x2255;
a1104<=x91 xor x498 xor x761 xor x1130 xor x1207 xor x2256;
a1105<=x92 xor x499 xor x762 xor x1131 xor x1208 xor x2257;
a1106<=x93 xor x500 xor x763 xor x1132 xor x1209 xor x2258;
a1107<=x94 xor x501 xor x764 xor x1133 xor x1210 xor x2259;
a1108<=x95 xor x502 xor x765 xor x1134 xor x1211 xor x2260;
a1109<=x96 xor x503 xor x766 xor x1135 xor x1212 xor x2261;
a1110<=x1 xor x504 xor x767 xor x1136 xor x1213 xor x2262;
a1111<=x2 xor x505 xor x768 xor x1137 xor x1214 xor x2263;
a1112<=x3 xor x506 xor x673 xor x1138 xor x1215 xor x2264;
a1113<=x4 xor x507 xor x674 xor x1139 xor x1216 xor x2265;
a1114<=x5 xor x508 xor x675 xor x1140 xor x1217 xor x2266;
a1115<=x6 xor x509 xor x676 xor x1141 xor x1218 xor x2267;
a1116<=x7 xor x510 xor x677 xor x1142 xor x1219 xor x2268;
a1117<=x8 xor x511 xor x678 xor x1143 xor x1220 xor x2269;
a1118<=x9 xor x512 xor x679 xor x1144 xor x1221 xor x2270;
a1119<=x10 xor x513 xor x680 xor x1145 xor x1222 xor x2271;
a1120<=x11 xor x514 xor x681 xor x1146 xor x1223 xor x2272;
a1121<=x12 xor x515 xor x682 xor x1147 xor x1224 xor x2273;
a1122<=x13 xor x516 xor x683 xor x1148 xor x1225 xor x2274;
a1123<=x14 xor x517 xor x684 xor x1149 xor x1226 xor x2275;
a1124<=x15 xor x518 xor x685 xor x1150 xor x1227 xor x2276;
a1125<=x16 xor x519 xor x686 xor x1151 xor x1228 xor x2277;
a1126<=x17 xor x520 xor x687 xor x1152 xor x1229 xor x2278;
a1127<=x18 xor x521 xor x688 xor x1057 xor x1230 xor x2279;
a1128<=x19 xor x522 xor x689 xor x1058 xor x1231 xor x2280;
a1129<=x20 xor x523 xor x690 xor x1059 xor x1232 xor x2281;
a1130<=x21 xor x524 xor x691 xor x1060 xor x1233 xor x2282;
a1131<=x22 xor x525 xor x692 xor x1061 xor x1234 xor x2283;
a1132<=x23 xor x526 xor x693 xor x1062 xor x1235 xor x2284;
a1133<=x24 xor x527 xor x694 xor x1063 xor x1236 xor x2285;
a1134<=x25 xor x528 xor x695 xor x1064 xor x1237 xor x2286;
a1135<=x26 xor x529 xor x696 xor x1065 xor x1238 xor x2287;
a1136<=x27 xor x530 xor x697 xor x1066 xor x1239 xor x2288;
a1137<=x28 xor x531 xor x698 xor x1067 xor x1240 xor x2289;
a1138<=x29 xor x532 xor x699 xor x1068 xor x1241 xor x2290;
a1139<=x30 xor x533 xor x700 xor x1069 xor x1242 xor x2291;
a1140<=x31 xor x534 xor x701 xor x1070 xor x1243 xor x2292;
a1141<=x32 xor x535 xor x702 xor x1071 xor x1244 xor x2293;
a1142<=x33 xor x536 xor x703 xor x1072 xor x1245 xor x2294;
a1143<=x34 xor x537 xor x704 xor x1073 xor x1246 xor x2295;
a1144<=x35 xor x538 xor x705 xor x1074 xor x1247 xor x2296;
a1145<=x36 xor x539 xor x706 xor x1075 xor x1248 xor x2297;
a1146<=x37 xor x540 xor x707 xor x1076 xor x1153 xor x2298;
a1147<=x38 xor x541 xor x708 xor x1077 xor x1154 xor x2299;
a1148<=x39 xor x542 xor x709 xor x1078 xor x1155 xor x2300;
a1149<=x40 xor x543 xor x710 xor x1079 xor x1156 xor x2301;
a1150<=x41 xor x544 xor x711 xor x1080 xor x1157 xor x2302;
a1151<=x42 xor x545 xor x712 xor x1081 xor x1158 xor x2303;
a1152<=x43 xor x546 xor x713 xor x1082 xor x1159 xor x2304;
Par<=a1 or a2 or a3 or a4 or a5 or a6 or a7 or a8 or a9 or a10 or a11 or a12 or a13 or a14 or a15 or a16 or a17 or a18 or a19 or a20 or a21 or a22 or a23 or a24 or a25 or a26 or a27 or a28 or a29 or a30 or a31 or a32 or a33 or a34 or a35 or a36 or a37 or a38 or a39 or a40 or a41 or a42 or a43 or a44 or a45 or a46 or a47 or a48 or a49 or a50 or a51 or a52 or a53 or a54 or a55 or a56 or a57 or a58 or a59 or a60 or a61 or a62 or a63 or a64 or a65 or a66 or a67 or a68 or a69 or a70 or a71 or a72 or a73 or a74 or a75 or a76 or a77 or a78 or a79 or a80 or a81 or a82 or a83 or a84 or a85 or a86 or a87 or a88 or a89 or a90 or a91 or a92 or a93 or a94 or a95 or a96 or a97 or a98 or a99 or a100 or a101 or a102 or a103 or a104 or a105 or a106 or a107 or a108 or a109 or a110 or a111 or a112 or a113 or a114 or a115 or a116 or a117 or a118 or a119 or a120 or a121 or a122 or a123 or a124 or a125 or a126 or a127 or a128 or a129 or a130 or a131 or a132 or a133 or a134 or a135 or a136 or a137 or a138 or a139 or a140 or a141 or a142 or a143 or a144 or a145 or a146 or a147 or a148 or a149 or a150 or a151 or a152 or a153 or a154 or a155 or a156 or a157 or a158 or a159 or a160 or a161 or a162 or a163 or a164 or a165 or a166 or a167 or a168 or a169 or a170 or a171 or a172 or a173 or a174 or a175 or a176 or a177 or a178 or a179 or a180 or a181 or a182 or a183 or a184 or a185 or a186 or a187 or a188 or a189 or a190 or a191 or a192 or a193 or a194 or a195 or a196 or a197 or a198 or a199 or a200 or a201 or a202 or a203 or a204 or a205 or a206 or a207 or a208 or a209 or a210 or a211 or a212 or a213 or a214 or a215 or a216 or a217 or a218 or a219 or a220 or a221 or a222 or a223 or a224 or a225 or a226 or a227 or a228 or a229 or a230 or a231 or a232 or a233 or a234 or a235 or a236 or a237 or a238 or a239 or a240 or a241 or a242 or a243 or a244 or a245 or a246 or a247 or a248 or a249 or a250 or a251 or a252 or a253 or a254 or a255 or a256 or a257 or a258 or a259 or a260 or a261 or a262 or a263 or a264 or a265 or a266 or a267 or a268 or a269 or a270 or a271 or a272 or a273 or a274 or a275 or a276 or a277 or a278 or a279 or a280 or a281 or a282 or a283 or a284 or a285 or a286 or a287 or a288 or a289 or a290 or a291 or a292 or a293 or a294 or a295 or a296 or a297 or a298 or a299 or a300 or a301 or a302 or a303 or a304 or a305 or a306 or a307 or a308 or a309 or a310 or a311 or a312 or a313 or a314 or a315 or a316 or a317 or a318 or a319 or a320 or a321 or a322 or a323 or a324 or a325 or a326 or a327 or a328 or a329 or a330 or a331 or a332 or a333 or a334 or a335 or a336 or a337 or a338 or a339 or a340 or a341 or a342 or a343 or a344 or a345 or a346 or a347 or a348 or a349 or a350 or a351 or a352 or a353 or a354 or a355 or a356 or a357 or a358 or a359 or a360 or a361 or a362 or a363 or a364 or a365 or a366 or a367 or a368 or a369 or a370 or a371 or a372 or a373 or a374 or a375 or a376 or a377 or a378 or a379 or a380 or a381 or a382 or a383 or a384 or a385 or a386 or a387 or a388 or a389 or a390 or a391 or a392 or a393 or a394 or a395 or a396 or a397 or a398 or a399 or a400 or a401 or a402 or a403 or a404 or a405 or a406 or a407 or a408 or a409 or a410 or a411 or a412 or a413 or a414 or a415 or a416 or a417 or a418 or a419 or a420 or a421 or a422 or a423 or a424 or a425 or a426 or a427 or a428 or a429 or a430 or a431 or a432 or a433 or a434 or a435 or a436 or a437 or a438 or a439 or a440 or a441 or a442 or a443 or a444 or a445 or a446 or a447 or a448 or a449 or a450 or a451 or a452 or a453 or a454 or a455 or a456 or a457 or a458 or a459 or a460 or a461 or a462 or a463 or a464 or a465 or a466 or a467 or a468 or a469 or a470 or a471 or a472 or a473 or a474 or a475 or a476 or a477 or a478 or a479 or a480 or a481 or a482 or a483 or a484 or a485 or a486 or a487 or a488 or a489 or a490 or a491 or a492 or a493 or a494 or a495 or a496 or a497 or a498 or a499 or a500 or a501 or a502 or a503 or a504 or a505 or a506 or a507 or a508 or a509 or a510 or a511 or a512 or a513 or a514 or a515 or a516 or a517 or a518 or a519 or a520 or a521 or a522 or a523 or a524 or a525 or a526 or a527 or a528 or a529 or a530 or a531 or a532 or a533 or a534 or a535 or a536 or a537 or a538 or a539 or a540 or a541 or a542 or a543 or a544 or a545 or a546 or a547 or a548 or a549 or a550 or a551 or a552 or a553 or a554 or a555 or a556 or a557 or a558 or a559 or a560 or a561 or a562 or a563 or a564 or a565 or a566 or a567 or a568 or a569 or a570 or a571 or a572 or a573 or a574 or a575 or a576 or a577 or a578 or a579 or a580 or a581 or a582 or a583 or a584 or a585 or a586 or a587 or a588 or a589 or a590 or a591 or a592 or a593 or a594 or a595 or a596 or a597 or a598 or a599 or a600 or a601 or a602 or a603 or a604 or a605 or a606 or a607 or a608 or a609 or a610 or a611 or a612 or a613 or a614 or a615 or a616 or a617 or a618 or a619 or a620 or a621 or a622 or a623 or a624 or a625 or a626 or a627 or a628 or a629 or a630 or a631 or a632 or a633 or a634 or a635 or a636 or a637 or a638 or a639 or a640 or a641 or a642 or a643 or a644 or a645 or a646 or a647 or a648 or a649 or a650 or a651 or a652 or a653 or a654 or a655 or a656 or a657 or a658 or a659 or a660 or a661 or a662 or a663 or a664 or a665 or a666 or a667 or a668 or a669 or a670 or a671 or a672 or a673 or a674 or a675 or a676 or a677 or a678 or a679 or a680 or a681 or a682 or a683 or a684 or a685 or a686 or a687 or a688 or a689 or a690 or a691 or a692 or a693 or a694 or a695 or a696 or a697 or a698 or a699 or a700 or a701 or a702 or a703 or a704 or a705 or a706 or a707 or a708 or a709 or a710 or a711 or a712 or a713 or a714 or a715 or a716 or a717 or a718 or a719 or a720 or a721 or a722 or a723 or a724 or a725 or a726 or a727 or a728 or a729 or a730 or a731 or a732 or a733 or a734 or a735 or a736 or a737 or a738 or a739 or a740 or a741 or a742 or a743 or a744 or a745 or a746 or a747 or a748 or a749 or a750 or a751 or a752 or a753 or a754 or a755 or a756 or a757 or a758 or a759 or a760 or a761 or a762 or a763 or a764 or a765 or a766 or a767 or a768 or a769 or a770 or a771 or a772 or a773 or a774 or a775 or a776 or a777 or a778 or a779 or a780 or a781 or a782 or a783 or a784 or a785 or a786 or a787 or a788 or a789 or a790 or a791 or a792 or a793 or a794 or a795 or a796 or a797 or a798 or a799 or a800 or a801 or a802 or a803 or a804 or a805 or a806 or a807 or a808 or a809 or a810 or a811 or a812 or a813 or a814 or a815 or a816 or a817 or a818 or a819 or a820 or a821 or a822 or a823 or a824 or a825 or a826 or a827 or a828 or a829 or a830 or a831 or a832 or a833 or a834 or a835 or a836 or a837 or a838 or a839 or a840 or a841 or a842 or a843 or a844 or a845 or a846 or a847 or a848 or a849 or a850 or a851 or a852 or a853 or a854 or a855 or a856 or a857 or a858 or a859 or a860 or a861 or a862 or a863 or a864 or a865 or a866 or a867 or a868 or a869 or a870 or a871 or a872 or a873 or a874 or a875 or a876 or a877 or a878 or a879 or a880 or a881 or a882 or a883 or a884 or a885 or a886 or a887 or a888 or a889 or a890 or a891 or a892 or a893 or a894 or a895 or a896 or a897 or a898 or a899 or a900 or a901 or a902 or a903 or a904 or a905 or a906 or a907 or a908 or a909 or a910 or a911 or a912 or a913 or a914 or a915 or a916 or a917 or a918 or a919 or a920 or a921 or a922 or a923 or a924 or a925 or a926 or a927 or a928 or a929 or a930 or a931 or a932 or a933 or a934 or a935 or a936 or a937 or a938 or a939 or a940 or a941 or a942 or a943 or a944 or a945 or a946 or a947 or a948 or a949 or a950 or a951 or a952 or a953 or a954 or a955 or a956 or a957 or a958 or a959 or a960 or a961 or a962 or a963 or a964 or a965 or a966 or a967 or a968 or a969 or a970 or a971 or a972 or a973 or a974 or a975 or a976 or a977 or a978 or a979 or a980 or a981 or a982 or a983 or a984 or a985 or a986 or a987 or a988 or a989 or a990 or a991 or a992 or a993 or a994 or a995 or a996 or a997 or a998 or a999 or a1000 or a1001 or a1002 or a1003 or a1004 or a1005 or a1006 or a1007 or a1008 or a1009 or a1010 or a1011 or a1012 or a1013 or a1014 or a1015 or a1016 or a1017 or a1018 or a1019 or a1020 or a1021 or a1022 or a1023 or a1024 or a1025 or a1026 or a1027 or a1028 or a1029 or a1030 or a1031 or a1032 or a1033 or a1034 or a1035 or a1036 or a1037 or a1038 or a1039 or a1040 or a1041 or a1042 or a1043 or a1044 or a1045 or a1046 or a1047 or a1048 or a1049 or a1050 or a1051 or a1052 or a1053 or a1054 or a1055 or a1056 or a1057 or a1058 or a1059 or a1060 or a1061 or a1062 or a1063 or a1064 or a1065 or a1066 or a1067 or a1068 or a1069 or a1070 or a1071 or a1072 or a1073 or a1074 or a1075 or a1076 or a1077 or a1078 or a1079 or a1080 or a1081 or a1082 or a1083 or a1084 or a1085 or a1086 or a1087 or a1088 or a1089 or a1090 or a1091 or a1092 or a1093 or a1094 or a1095 or a1096 or a1097 or a1098 or a1099 or a1100 or a1101 or a1102 or a1103 or a1104 or a1105 or a1106 or a1107 or a1108 or a1109 or a1110 or a1111 or a1112 or a1113 or a1114 or a1115 or a1116 or a1117 or a1118 or a1119 or a1120 or a1121 or a1122 or a1123 or a1124 or a1125 or a1126 or a1127 or a1128 or a1129 or a1130 or a1131 or a1132 or a1133 or a1134 or a1135 or a1136 or a1137 or a1138 or a1139 or a1140 or a1141 or a1142 or a1143 or a1144 or a1145 or a1146 or a1147 or a1148 or a1149 or a1150 or a1151 or a1152;
 
process(clk,start_pa,rst,count,itmax)
begin
if(rst='1') then
count<="00000";
elsif(rising_edge(clk) and start_pa='1')then
count<=count+1;
else 
count<=count;
end if;
end process;
nbr_iter<=std_logic_vector(count);
end_decision<='1' when count>=itmax or Par='0' else '0';
end;