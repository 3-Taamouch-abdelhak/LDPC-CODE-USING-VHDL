LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY decoder IS PORT(
     clock,reset,start_decoder   :in std_logic;
     iter_Mx          :in    std_logic_vector(4 downto 0);
     L1              :in std_logic_vector(8 DOWNTO 0);
     L2              :in std_logic_vector(8 DOWNTO 0);
     L3              :in std_logic_vector(8 DOWNTO 0);
     L4              :in std_logic_vector(8 DOWNTO 0);
     L5              :in std_logic_vector(8 DOWNTO 0);
     L6              :in std_logic_vector(8 DOWNTO 0);
     L7              :in std_logic_vector(8 DOWNTO 0);
     L8              :in std_logic_vector(8 DOWNTO 0);
     L9              :in std_logic_vector(8 DOWNTO 0);
     L10              :in std_logic_vector(8 DOWNTO 0);
     L11              :in std_logic_vector(8 DOWNTO 0);
     L12              :in std_logic_vector(8 DOWNTO 0);
     L13              :in std_logic_vector(8 DOWNTO 0);
     L14              :in std_logic_vector(8 DOWNTO 0);
     L15              :in std_logic_vector(8 DOWNTO 0);
     L16              :in std_logic_vector(8 DOWNTO 0);
     L17              :in std_logic_vector(8 DOWNTO 0);
     L18              :in std_logic_vector(8 DOWNTO 0);
     L19              :in std_logic_vector(8 DOWNTO 0);
     L20              :in std_logic_vector(8 DOWNTO 0);
     L21              :in std_logic_vector(8 DOWNTO 0);
     L22              :in std_logic_vector(8 DOWNTO 0);
     L23              :in std_logic_vector(8 DOWNTO 0);
     L24              :in std_logic_vector(8 DOWNTO 0);
     L25              :in std_logic_vector(8 DOWNTO 0);
     L26              :in std_logic_vector(8 DOWNTO 0);
     L27              :in std_logic_vector(8 DOWNTO 0);
     L28              :in std_logic_vector(8 DOWNTO 0);
     L29              :in std_logic_vector(8 DOWNTO 0);
     L30              :in std_logic_vector(8 DOWNTO 0);
     L31              :in std_logic_vector(8 DOWNTO 0);
     L32              :in std_logic_vector(8 DOWNTO 0);
     L33              :in std_logic_vector(8 DOWNTO 0);
     L34              :in std_logic_vector(8 DOWNTO 0);
     L35              :in std_logic_vector(8 DOWNTO 0);
     L36              :in std_logic_vector(8 DOWNTO 0);
     L37              :in std_logic_vector(8 DOWNTO 0);
     L38              :in std_logic_vector(8 DOWNTO 0);
     L39              :in std_logic_vector(8 DOWNTO 0);
     L40              :in std_logic_vector(8 DOWNTO 0);
     L41              :in std_logic_vector(8 DOWNTO 0);
     L42              :in std_logic_vector(8 DOWNTO 0);
     L43              :in std_logic_vector(8 DOWNTO 0);
     L44              :in std_logic_vector(8 DOWNTO 0);
     L45              :in std_logic_vector(8 DOWNTO 0);
     L46              :in std_logic_vector(8 DOWNTO 0);
     L47              :in std_logic_vector(8 DOWNTO 0);
     L48              :in std_logic_vector(8 DOWNTO 0);
     L49              :in std_logic_vector(8 DOWNTO 0);
     L50              :in std_logic_vector(8 DOWNTO 0);
     L51              :in std_logic_vector(8 DOWNTO 0);
     L52              :in std_logic_vector(8 DOWNTO 0);
     L53              :in std_logic_vector(8 DOWNTO 0);
     L54              :in std_logic_vector(8 DOWNTO 0);
     L55              :in std_logic_vector(8 DOWNTO 0);
     L56              :in std_logic_vector(8 DOWNTO 0);
     L57              :in std_logic_vector(8 DOWNTO 0);
     L58              :in std_logic_vector(8 DOWNTO 0);
     L59              :in std_logic_vector(8 DOWNTO 0);
     L60              :in std_logic_vector(8 DOWNTO 0);
     L61              :in std_logic_vector(8 DOWNTO 0);
     L62              :in std_logic_vector(8 DOWNTO 0);
     L63              :in std_logic_vector(8 DOWNTO 0);
     L64              :in std_logic_vector(8 DOWNTO 0);
     L65              :in std_logic_vector(8 DOWNTO 0);
     L66              :in std_logic_vector(8 DOWNTO 0);
     L67              :in std_logic_vector(8 DOWNTO 0);
     L68              :in std_logic_vector(8 DOWNTO 0);
     L69              :in std_logic_vector(8 DOWNTO 0);
     L70              :in std_logic_vector(8 DOWNTO 0);
     L71              :in std_logic_vector(8 DOWNTO 0);
     L72              :in std_logic_vector(8 DOWNTO 0);
     L73              :in std_logic_vector(8 DOWNTO 0);
     L74              :in std_logic_vector(8 DOWNTO 0);
     L75              :in std_logic_vector(8 DOWNTO 0);
     L76              :in std_logic_vector(8 DOWNTO 0);
     L77              :in std_logic_vector(8 DOWNTO 0);
     L78              :in std_logic_vector(8 DOWNTO 0);
     L79              :in std_logic_vector(8 DOWNTO 0);
     L80              :in std_logic_vector(8 DOWNTO 0);
     L81              :in std_logic_vector(8 DOWNTO 0);
     L82              :in std_logic_vector(8 DOWNTO 0);
     L83              :in std_logic_vector(8 DOWNTO 0);
     L84              :in std_logic_vector(8 DOWNTO 0);
     L85              :in std_logic_vector(8 DOWNTO 0);
     L86              :in std_logic_vector(8 DOWNTO 0);
     L87              :in std_logic_vector(8 DOWNTO 0);
     L88              :in std_logic_vector(8 DOWNTO 0);
     L89              :in std_logic_vector(8 DOWNTO 0);
     L90              :in std_logic_vector(8 DOWNTO 0);
     L91              :in std_logic_vector(8 DOWNTO 0);
     L92              :in std_logic_vector(8 DOWNTO 0);
     L93              :in std_logic_vector(8 DOWNTO 0);
     L94              :in std_logic_vector(8 DOWNTO 0);
     L95              :in std_logic_vector(8 DOWNTO 0);
     L96              :in std_logic_vector(8 DOWNTO 0);
     L97              :in std_logic_vector(8 DOWNTO 0);
     L98              :in std_logic_vector(8 DOWNTO 0);
     L99              :in std_logic_vector(8 DOWNTO 0);
     L100              :in std_logic_vector(8 DOWNTO 0);
     L101              :in std_logic_vector(8 DOWNTO 0);
     L102              :in std_logic_vector(8 DOWNTO 0);
     L103              :in std_logic_vector(8 DOWNTO 0);
     L104              :in std_logic_vector(8 DOWNTO 0);
     L105              :in std_logic_vector(8 DOWNTO 0);
     L106              :in std_logic_vector(8 DOWNTO 0);
     L107              :in std_logic_vector(8 DOWNTO 0);
     L108              :in std_logic_vector(8 DOWNTO 0);
     L109              :in std_logic_vector(8 DOWNTO 0);
     L110              :in std_logic_vector(8 DOWNTO 0);
     L111              :in std_logic_vector(8 DOWNTO 0);
     L112              :in std_logic_vector(8 DOWNTO 0);
     L113              :in std_logic_vector(8 DOWNTO 0);
     L114              :in std_logic_vector(8 DOWNTO 0);
     L115              :in std_logic_vector(8 DOWNTO 0);
     L116              :in std_logic_vector(8 DOWNTO 0);
     L117              :in std_logic_vector(8 DOWNTO 0);
     L118              :in std_logic_vector(8 DOWNTO 0);
     L119              :in std_logic_vector(8 DOWNTO 0);
     L120              :in std_logic_vector(8 DOWNTO 0);
     L121              :in std_logic_vector(8 DOWNTO 0);
     L122              :in std_logic_vector(8 DOWNTO 0);
     L123              :in std_logic_vector(8 DOWNTO 0);
     L124              :in std_logic_vector(8 DOWNTO 0);
     L125              :in std_logic_vector(8 DOWNTO 0);
     L126              :in std_logic_vector(8 DOWNTO 0);
     L127              :in std_logic_vector(8 DOWNTO 0);
     L128              :in std_logic_vector(8 DOWNTO 0);
     L129              :in std_logic_vector(8 DOWNTO 0);
     L130              :in std_logic_vector(8 DOWNTO 0);
     L131              :in std_logic_vector(8 DOWNTO 0);
     L132              :in std_logic_vector(8 DOWNTO 0);
     L133              :in std_logic_vector(8 DOWNTO 0);
     L134              :in std_logic_vector(8 DOWNTO 0);
     L135              :in std_logic_vector(8 DOWNTO 0);
     L136              :in std_logic_vector(8 DOWNTO 0);
     L137              :in std_logic_vector(8 DOWNTO 0);
     L138              :in std_logic_vector(8 DOWNTO 0);
     L139              :in std_logic_vector(8 DOWNTO 0);
     L140              :in std_logic_vector(8 DOWNTO 0);
     L141              :in std_logic_vector(8 DOWNTO 0);
     L142              :in std_logic_vector(8 DOWNTO 0);
     L143              :in std_logic_vector(8 DOWNTO 0);
     L144              :in std_logic_vector(8 DOWNTO 0);
     L145              :in std_logic_vector(8 DOWNTO 0);
     L146              :in std_logic_vector(8 DOWNTO 0);
     L147              :in std_logic_vector(8 DOWNTO 0);
     L148              :in std_logic_vector(8 DOWNTO 0);
     L149              :in std_logic_vector(8 DOWNTO 0);
     L150              :in std_logic_vector(8 DOWNTO 0);
     L151              :in std_logic_vector(8 DOWNTO 0);
     L152              :in std_logic_vector(8 DOWNTO 0);
     L153              :in std_logic_vector(8 DOWNTO 0);
     L154              :in std_logic_vector(8 DOWNTO 0);
     L155              :in std_logic_vector(8 DOWNTO 0);
     L156              :in std_logic_vector(8 DOWNTO 0);
     L157              :in std_logic_vector(8 DOWNTO 0);
     L158              :in std_logic_vector(8 DOWNTO 0);
     L159              :in std_logic_vector(8 DOWNTO 0);
     L160              :in std_logic_vector(8 DOWNTO 0);
     L161              :in std_logic_vector(8 DOWNTO 0);
     L162              :in std_logic_vector(8 DOWNTO 0);
     L163              :in std_logic_vector(8 DOWNTO 0);
     L164              :in std_logic_vector(8 DOWNTO 0);
     L165              :in std_logic_vector(8 DOWNTO 0);
     L166              :in std_logic_vector(8 DOWNTO 0);
     L167              :in std_logic_vector(8 DOWNTO 0);
     L168              :in std_logic_vector(8 DOWNTO 0);
     L169              :in std_logic_vector(8 DOWNTO 0);
     L170              :in std_logic_vector(8 DOWNTO 0);
     L171              :in std_logic_vector(8 DOWNTO 0);
     L172              :in std_logic_vector(8 DOWNTO 0);
     L173              :in std_logic_vector(8 DOWNTO 0);
     L174              :in std_logic_vector(8 DOWNTO 0);
     L175              :in std_logic_vector(8 DOWNTO 0);
     L176              :in std_logic_vector(8 DOWNTO 0);
     L177              :in std_logic_vector(8 DOWNTO 0);
     L178              :in std_logic_vector(8 DOWNTO 0);
     L179              :in std_logic_vector(8 DOWNTO 0);
     L180              :in std_logic_vector(8 DOWNTO 0);
     L181              :in std_logic_vector(8 DOWNTO 0);
     L182              :in std_logic_vector(8 DOWNTO 0);
     L183              :in std_logic_vector(8 DOWNTO 0);
     L184              :in std_logic_vector(8 DOWNTO 0);
     L185              :in std_logic_vector(8 DOWNTO 0);
     L186              :in std_logic_vector(8 DOWNTO 0);
     L187              :in std_logic_vector(8 DOWNTO 0);
     L188              :in std_logic_vector(8 DOWNTO 0);
     L189              :in std_logic_vector(8 DOWNTO 0);
     L190              :in std_logic_vector(8 DOWNTO 0);
     L191              :in std_logic_vector(8 DOWNTO 0);
     L192              :in std_logic_vector(8 DOWNTO 0);
     L193              :in std_logic_vector(8 DOWNTO 0);
     L194              :in std_logic_vector(8 DOWNTO 0);
     L195              :in std_logic_vector(8 DOWNTO 0);
     L196              :in std_logic_vector(8 DOWNTO 0);
     L197              :in std_logic_vector(8 DOWNTO 0);
     L198              :in std_logic_vector(8 DOWNTO 0);
     L199              :in std_logic_vector(8 DOWNTO 0);
     L200              :in std_logic_vector(8 DOWNTO 0);
     L201              :in std_logic_vector(8 DOWNTO 0);
     L202              :in std_logic_vector(8 DOWNTO 0);
     L203              :in std_logic_vector(8 DOWNTO 0);
     L204              :in std_logic_vector(8 DOWNTO 0);
     L205              :in std_logic_vector(8 DOWNTO 0);
     L206              :in std_logic_vector(8 DOWNTO 0);
     L207              :in std_logic_vector(8 DOWNTO 0);
     L208              :in std_logic_vector(8 DOWNTO 0);
     L209              :in std_logic_vector(8 DOWNTO 0);
     L210              :in std_logic_vector(8 DOWNTO 0);
     L211              :in std_logic_vector(8 DOWNTO 0);
     L212              :in std_logic_vector(8 DOWNTO 0);
     L213              :in std_logic_vector(8 DOWNTO 0);
     L214              :in std_logic_vector(8 DOWNTO 0);
     L215              :in std_logic_vector(8 DOWNTO 0);
     L216              :in std_logic_vector(8 DOWNTO 0);
     L217              :in std_logic_vector(8 DOWNTO 0);
     L218              :in std_logic_vector(8 DOWNTO 0);
     L219              :in std_logic_vector(8 DOWNTO 0);
     L220              :in std_logic_vector(8 DOWNTO 0);
     L221              :in std_logic_vector(8 DOWNTO 0);
     L222              :in std_logic_vector(8 DOWNTO 0);
     L223              :in std_logic_vector(8 DOWNTO 0);
     L224              :in std_logic_vector(8 DOWNTO 0);
     L225              :in std_logic_vector(8 DOWNTO 0);
     L226              :in std_logic_vector(8 DOWNTO 0);
     L227              :in std_logic_vector(8 DOWNTO 0);
     L228              :in std_logic_vector(8 DOWNTO 0);
     L229              :in std_logic_vector(8 DOWNTO 0);
     L230              :in std_logic_vector(8 DOWNTO 0);
     L231              :in std_logic_vector(8 DOWNTO 0);
     L232              :in std_logic_vector(8 DOWNTO 0);
     L233              :in std_logic_vector(8 DOWNTO 0);
     L234              :in std_logic_vector(8 DOWNTO 0);
     L235              :in std_logic_vector(8 DOWNTO 0);
     L236              :in std_logic_vector(8 DOWNTO 0);
     L237              :in std_logic_vector(8 DOWNTO 0);
     L238              :in std_logic_vector(8 DOWNTO 0);
     L239              :in std_logic_vector(8 DOWNTO 0);
     L240              :in std_logic_vector(8 DOWNTO 0);
     L241              :in std_logic_vector(8 DOWNTO 0);
     L242              :in std_logic_vector(8 DOWNTO 0);
     L243              :in std_logic_vector(8 DOWNTO 0);
     L244              :in std_logic_vector(8 DOWNTO 0);
     L245              :in std_logic_vector(8 DOWNTO 0);
     L246              :in std_logic_vector(8 DOWNTO 0);
     L247              :in std_logic_vector(8 DOWNTO 0);
     L248              :in std_logic_vector(8 DOWNTO 0);
     L249              :in std_logic_vector(8 DOWNTO 0);
     L250              :in std_logic_vector(8 DOWNTO 0);
     L251              :in std_logic_vector(8 DOWNTO 0);
     L252              :in std_logic_vector(8 DOWNTO 0);
     L253              :in std_logic_vector(8 DOWNTO 0);
     L254              :in std_logic_vector(8 DOWNTO 0);
     L255              :in std_logic_vector(8 DOWNTO 0);
     L256              :in std_logic_vector(8 DOWNTO 0);
     L257              :in std_logic_vector(8 DOWNTO 0);
     L258              :in std_logic_vector(8 DOWNTO 0);
     L259              :in std_logic_vector(8 DOWNTO 0);
     L260              :in std_logic_vector(8 DOWNTO 0);
     L261              :in std_logic_vector(8 DOWNTO 0);
     L262              :in std_logic_vector(8 DOWNTO 0);
     L263              :in std_logic_vector(8 DOWNTO 0);
     L264              :in std_logic_vector(8 DOWNTO 0);
     L265              :in std_logic_vector(8 DOWNTO 0);
     L266              :in std_logic_vector(8 DOWNTO 0);
     L267              :in std_logic_vector(8 DOWNTO 0);
     L268              :in std_logic_vector(8 DOWNTO 0);
     L269              :in std_logic_vector(8 DOWNTO 0);
     L270              :in std_logic_vector(8 DOWNTO 0);
     L271              :in std_logic_vector(8 DOWNTO 0);
     L272              :in std_logic_vector(8 DOWNTO 0);
     L273              :in std_logic_vector(8 DOWNTO 0);
     L274              :in std_logic_vector(8 DOWNTO 0);
     L275              :in std_logic_vector(8 DOWNTO 0);
     L276              :in std_logic_vector(8 DOWNTO 0);
     L277              :in std_logic_vector(8 DOWNTO 0);
     L278              :in std_logic_vector(8 DOWNTO 0);
     L279              :in std_logic_vector(8 DOWNTO 0);
     L280              :in std_logic_vector(8 DOWNTO 0);
     L281              :in std_logic_vector(8 DOWNTO 0);
     L282              :in std_logic_vector(8 DOWNTO 0);
     L283              :in std_logic_vector(8 DOWNTO 0);
     L284              :in std_logic_vector(8 DOWNTO 0);
     L285              :in std_logic_vector(8 DOWNTO 0);
     L286              :in std_logic_vector(8 DOWNTO 0);
     L287              :in std_logic_vector(8 DOWNTO 0);
     L288              :in std_logic_vector(8 DOWNTO 0);
     L289              :in std_logic_vector(8 DOWNTO 0);
     L290              :in std_logic_vector(8 DOWNTO 0);
     L291              :in std_logic_vector(8 DOWNTO 0);
     L292              :in std_logic_vector(8 DOWNTO 0);
     L293              :in std_logic_vector(8 DOWNTO 0);
     L294              :in std_logic_vector(8 DOWNTO 0);
     L295              :in std_logic_vector(8 DOWNTO 0);
     L296              :in std_logic_vector(8 DOWNTO 0);
     L297              :in std_logic_vector(8 DOWNTO 0);
     L298              :in std_logic_vector(8 DOWNTO 0);
     L299              :in std_logic_vector(8 DOWNTO 0);
     L300              :in std_logic_vector(8 DOWNTO 0);
     L301              :in std_logic_vector(8 DOWNTO 0);
     L302              :in std_logic_vector(8 DOWNTO 0);
     L303              :in std_logic_vector(8 DOWNTO 0);
     L304              :in std_logic_vector(8 DOWNTO 0);
     L305              :in std_logic_vector(8 DOWNTO 0);
     L306              :in std_logic_vector(8 DOWNTO 0);
     L307              :in std_logic_vector(8 DOWNTO 0);
     L308              :in std_logic_vector(8 DOWNTO 0);
     L309              :in std_logic_vector(8 DOWNTO 0);
     L310              :in std_logic_vector(8 DOWNTO 0);
     L311              :in std_logic_vector(8 DOWNTO 0);
     L312              :in std_logic_vector(8 DOWNTO 0);
     L313              :in std_logic_vector(8 DOWNTO 0);
     L314              :in std_logic_vector(8 DOWNTO 0);
     L315              :in std_logic_vector(8 DOWNTO 0);
     L316              :in std_logic_vector(8 DOWNTO 0);
     L317              :in std_logic_vector(8 DOWNTO 0);
     L318              :in std_logic_vector(8 DOWNTO 0);
     L319              :in std_logic_vector(8 DOWNTO 0);
     L320              :in std_logic_vector(8 DOWNTO 0);
     L321              :in std_logic_vector(8 DOWNTO 0);
     L322              :in std_logic_vector(8 DOWNTO 0);
     L323              :in std_logic_vector(8 DOWNTO 0);
     L324              :in std_logic_vector(8 DOWNTO 0);
     L325              :in std_logic_vector(8 DOWNTO 0);
     L326              :in std_logic_vector(8 DOWNTO 0);
     L327              :in std_logic_vector(8 DOWNTO 0);
     L328              :in std_logic_vector(8 DOWNTO 0);
     L329              :in std_logic_vector(8 DOWNTO 0);
     L330              :in std_logic_vector(8 DOWNTO 0);
     L331              :in std_logic_vector(8 DOWNTO 0);
     L332              :in std_logic_vector(8 DOWNTO 0);
     L333              :in std_logic_vector(8 DOWNTO 0);
     L334              :in std_logic_vector(8 DOWNTO 0);
     L335              :in std_logic_vector(8 DOWNTO 0);
     L336              :in std_logic_vector(8 DOWNTO 0);
     L337              :in std_logic_vector(8 DOWNTO 0);
     L338              :in std_logic_vector(8 DOWNTO 0);
     L339              :in std_logic_vector(8 DOWNTO 0);
     L340              :in std_logic_vector(8 DOWNTO 0);
     L341              :in std_logic_vector(8 DOWNTO 0);
     L342              :in std_logic_vector(8 DOWNTO 0);
     L343              :in std_logic_vector(8 DOWNTO 0);
     L344              :in std_logic_vector(8 DOWNTO 0);
     L345              :in std_logic_vector(8 DOWNTO 0);
     L346              :in std_logic_vector(8 DOWNTO 0);
     L347              :in std_logic_vector(8 DOWNTO 0);
     L348              :in std_logic_vector(8 DOWNTO 0);
     L349              :in std_logic_vector(8 DOWNTO 0);
     L350              :in std_logic_vector(8 DOWNTO 0);
     L351              :in std_logic_vector(8 DOWNTO 0);
     L352              :in std_logic_vector(8 DOWNTO 0);
     L353              :in std_logic_vector(8 DOWNTO 0);
     L354              :in std_logic_vector(8 DOWNTO 0);
     L355              :in std_logic_vector(8 DOWNTO 0);
     L356              :in std_logic_vector(8 DOWNTO 0);
     L357              :in std_logic_vector(8 DOWNTO 0);
     L358              :in std_logic_vector(8 DOWNTO 0);
     L359              :in std_logic_vector(8 DOWNTO 0);
     L360              :in std_logic_vector(8 DOWNTO 0);
     L361              :in std_logic_vector(8 DOWNTO 0);
     L362              :in std_logic_vector(8 DOWNTO 0);
     L363              :in std_logic_vector(8 DOWNTO 0);
     L364              :in std_logic_vector(8 DOWNTO 0);
     L365              :in std_logic_vector(8 DOWNTO 0);
     L366              :in std_logic_vector(8 DOWNTO 0);
     L367              :in std_logic_vector(8 DOWNTO 0);
     L368              :in std_logic_vector(8 DOWNTO 0);
     L369              :in std_logic_vector(8 DOWNTO 0);
     L370              :in std_logic_vector(8 DOWNTO 0);
     L371              :in std_logic_vector(8 DOWNTO 0);
     L372              :in std_logic_vector(8 DOWNTO 0);
     L373              :in std_logic_vector(8 DOWNTO 0);
     L374              :in std_logic_vector(8 DOWNTO 0);
     L375              :in std_logic_vector(8 DOWNTO 0);
     L376              :in std_logic_vector(8 DOWNTO 0);
     L377              :in std_logic_vector(8 DOWNTO 0);
     L378              :in std_logic_vector(8 DOWNTO 0);
     L379              :in std_logic_vector(8 DOWNTO 0);
     L380              :in std_logic_vector(8 DOWNTO 0);
     L381              :in std_logic_vector(8 DOWNTO 0);
     L382              :in std_logic_vector(8 DOWNTO 0);
     L383              :in std_logic_vector(8 DOWNTO 0);
     L384              :in std_logic_vector(8 DOWNTO 0);
     L385              :in std_logic_vector(8 DOWNTO 0);
     L386              :in std_logic_vector(8 DOWNTO 0);
     L387              :in std_logic_vector(8 DOWNTO 0);
     L388              :in std_logic_vector(8 DOWNTO 0);
     L389              :in std_logic_vector(8 DOWNTO 0);
     L390              :in std_logic_vector(8 DOWNTO 0);
     L391              :in std_logic_vector(8 DOWNTO 0);
     L392              :in std_logic_vector(8 DOWNTO 0);
     L393              :in std_logic_vector(8 DOWNTO 0);
     L394              :in std_logic_vector(8 DOWNTO 0);
     L395              :in std_logic_vector(8 DOWNTO 0);
     L396              :in std_logic_vector(8 DOWNTO 0);
     L397              :in std_logic_vector(8 DOWNTO 0);
     L398              :in std_logic_vector(8 DOWNTO 0);
     L399              :in std_logic_vector(8 DOWNTO 0);
     L400              :in std_logic_vector(8 DOWNTO 0);
     L401              :in std_logic_vector(8 DOWNTO 0);
     L402              :in std_logic_vector(8 DOWNTO 0);
     L403              :in std_logic_vector(8 DOWNTO 0);
     L404              :in std_logic_vector(8 DOWNTO 0);
     L405              :in std_logic_vector(8 DOWNTO 0);
     L406              :in std_logic_vector(8 DOWNTO 0);
     L407              :in std_logic_vector(8 DOWNTO 0);
     L408              :in std_logic_vector(8 DOWNTO 0);
     L409              :in std_logic_vector(8 DOWNTO 0);
     L410              :in std_logic_vector(8 DOWNTO 0);
     L411              :in std_logic_vector(8 DOWNTO 0);
     L412              :in std_logic_vector(8 DOWNTO 0);
     L413              :in std_logic_vector(8 DOWNTO 0);
     L414              :in std_logic_vector(8 DOWNTO 0);
     L415              :in std_logic_vector(8 DOWNTO 0);
     L416              :in std_logic_vector(8 DOWNTO 0);
     L417              :in std_logic_vector(8 DOWNTO 0);
     L418              :in std_logic_vector(8 DOWNTO 0);
     L419              :in std_logic_vector(8 DOWNTO 0);
     L420              :in std_logic_vector(8 DOWNTO 0);
     L421              :in std_logic_vector(8 DOWNTO 0);
     L422              :in std_logic_vector(8 DOWNTO 0);
     L423              :in std_logic_vector(8 DOWNTO 0);
     L424              :in std_logic_vector(8 DOWNTO 0);
     L425              :in std_logic_vector(8 DOWNTO 0);
     L426              :in std_logic_vector(8 DOWNTO 0);
     L427              :in std_logic_vector(8 DOWNTO 0);
     L428              :in std_logic_vector(8 DOWNTO 0);
     L429              :in std_logic_vector(8 DOWNTO 0);
     L430              :in std_logic_vector(8 DOWNTO 0);
     L431              :in std_logic_vector(8 DOWNTO 0);
     L432              :in std_logic_vector(8 DOWNTO 0);
     L433              :in std_logic_vector(8 DOWNTO 0);
     L434              :in std_logic_vector(8 DOWNTO 0);
     L435              :in std_logic_vector(8 DOWNTO 0);
     L436              :in std_logic_vector(8 DOWNTO 0);
     L437              :in std_logic_vector(8 DOWNTO 0);
     L438              :in std_logic_vector(8 DOWNTO 0);
     L439              :in std_logic_vector(8 DOWNTO 0);
     L440              :in std_logic_vector(8 DOWNTO 0);
     L441              :in std_logic_vector(8 DOWNTO 0);
     L442              :in std_logic_vector(8 DOWNTO 0);
     L443              :in std_logic_vector(8 DOWNTO 0);
     L444              :in std_logic_vector(8 DOWNTO 0);
     L445              :in std_logic_vector(8 DOWNTO 0);
     L446              :in std_logic_vector(8 DOWNTO 0);
     L447              :in std_logic_vector(8 DOWNTO 0);
     L448              :in std_logic_vector(8 DOWNTO 0);
     L449              :in std_logic_vector(8 DOWNTO 0);
     L450              :in std_logic_vector(8 DOWNTO 0);
     L451              :in std_logic_vector(8 DOWNTO 0);
     L452              :in std_logic_vector(8 DOWNTO 0);
     L453              :in std_logic_vector(8 DOWNTO 0);
     L454              :in std_logic_vector(8 DOWNTO 0);
     L455              :in std_logic_vector(8 DOWNTO 0);
     L456              :in std_logic_vector(8 DOWNTO 0);
     L457              :in std_logic_vector(8 DOWNTO 0);
     L458              :in std_logic_vector(8 DOWNTO 0);
     L459              :in std_logic_vector(8 DOWNTO 0);
     L460              :in std_logic_vector(8 DOWNTO 0);
     L461              :in std_logic_vector(8 DOWNTO 0);
     L462              :in std_logic_vector(8 DOWNTO 0);
     L463              :in std_logic_vector(8 DOWNTO 0);
     L464              :in std_logic_vector(8 DOWNTO 0);
     L465              :in std_logic_vector(8 DOWNTO 0);
     L466              :in std_logic_vector(8 DOWNTO 0);
     L467              :in std_logic_vector(8 DOWNTO 0);
     L468              :in std_logic_vector(8 DOWNTO 0);
     L469              :in std_logic_vector(8 DOWNTO 0);
     L470              :in std_logic_vector(8 DOWNTO 0);
     L471              :in std_logic_vector(8 DOWNTO 0);
     L472              :in std_logic_vector(8 DOWNTO 0);
     L473              :in std_logic_vector(8 DOWNTO 0);
     L474              :in std_logic_vector(8 DOWNTO 0);
     L475              :in std_logic_vector(8 DOWNTO 0);
     L476              :in std_logic_vector(8 DOWNTO 0);
     L477              :in std_logic_vector(8 DOWNTO 0);
     L478              :in std_logic_vector(8 DOWNTO 0);
     L479              :in std_logic_vector(8 DOWNTO 0);
     L480              :in std_logic_vector(8 DOWNTO 0);
     L481              :in std_logic_vector(8 DOWNTO 0);
     L482              :in std_logic_vector(8 DOWNTO 0);
     L483              :in std_logic_vector(8 DOWNTO 0);
     L484              :in std_logic_vector(8 DOWNTO 0);
     L485              :in std_logic_vector(8 DOWNTO 0);
     L486              :in std_logic_vector(8 DOWNTO 0);
     L487              :in std_logic_vector(8 DOWNTO 0);
     L488              :in std_logic_vector(8 DOWNTO 0);
     L489              :in std_logic_vector(8 DOWNTO 0);
     L490              :in std_logic_vector(8 DOWNTO 0);
     L491              :in std_logic_vector(8 DOWNTO 0);
     L492              :in std_logic_vector(8 DOWNTO 0);
     L493              :in std_logic_vector(8 DOWNTO 0);
     L494              :in std_logic_vector(8 DOWNTO 0);
     L495              :in std_logic_vector(8 DOWNTO 0);
     L496              :in std_logic_vector(8 DOWNTO 0);
     L497              :in std_logic_vector(8 DOWNTO 0);
     L498              :in std_logic_vector(8 DOWNTO 0);
     L499              :in std_logic_vector(8 DOWNTO 0);
     L500              :in std_logic_vector(8 DOWNTO 0);
     L501              :in std_logic_vector(8 DOWNTO 0);
     L502              :in std_logic_vector(8 DOWNTO 0);
     L503              :in std_logic_vector(8 DOWNTO 0);
     L504              :in std_logic_vector(8 DOWNTO 0);
     L505              :in std_logic_vector(8 DOWNTO 0);
     L506              :in std_logic_vector(8 DOWNTO 0);
     L507              :in std_logic_vector(8 DOWNTO 0);
     L508              :in std_logic_vector(8 DOWNTO 0);
     L509              :in std_logic_vector(8 DOWNTO 0);
     L510              :in std_logic_vector(8 DOWNTO 0);
     L511              :in std_logic_vector(8 DOWNTO 0);
     L512              :in std_logic_vector(8 DOWNTO 0);
     L513              :in std_logic_vector(8 DOWNTO 0);
     L514              :in std_logic_vector(8 DOWNTO 0);
     L515              :in std_logic_vector(8 DOWNTO 0);
     L516              :in std_logic_vector(8 DOWNTO 0);
     L517              :in std_logic_vector(8 DOWNTO 0);
     L518              :in std_logic_vector(8 DOWNTO 0);
     L519              :in std_logic_vector(8 DOWNTO 0);
     L520              :in std_logic_vector(8 DOWNTO 0);
     L521              :in std_logic_vector(8 DOWNTO 0);
     L522              :in std_logic_vector(8 DOWNTO 0);
     L523              :in std_logic_vector(8 DOWNTO 0);
     L524              :in std_logic_vector(8 DOWNTO 0);
     L525              :in std_logic_vector(8 DOWNTO 0);
     L526              :in std_logic_vector(8 DOWNTO 0);
     L527              :in std_logic_vector(8 DOWNTO 0);
     L528              :in std_logic_vector(8 DOWNTO 0);
     L529              :in std_logic_vector(8 DOWNTO 0);
     L530              :in std_logic_vector(8 DOWNTO 0);
     L531              :in std_logic_vector(8 DOWNTO 0);
     L532              :in std_logic_vector(8 DOWNTO 0);
     L533              :in std_logic_vector(8 DOWNTO 0);
     L534              :in std_logic_vector(8 DOWNTO 0);
     L535              :in std_logic_vector(8 DOWNTO 0);
     L536              :in std_logic_vector(8 DOWNTO 0);
     L537              :in std_logic_vector(8 DOWNTO 0);
     L538              :in std_logic_vector(8 DOWNTO 0);
     L539              :in std_logic_vector(8 DOWNTO 0);
     L540              :in std_logic_vector(8 DOWNTO 0);
     L541              :in std_logic_vector(8 DOWNTO 0);
     L542              :in std_logic_vector(8 DOWNTO 0);
     L543              :in std_logic_vector(8 DOWNTO 0);
     L544              :in std_logic_vector(8 DOWNTO 0);
     L545              :in std_logic_vector(8 DOWNTO 0);
     L546              :in std_logic_vector(8 DOWNTO 0);
     L547              :in std_logic_vector(8 DOWNTO 0);
     L548              :in std_logic_vector(8 DOWNTO 0);
     L549              :in std_logic_vector(8 DOWNTO 0);
     L550              :in std_logic_vector(8 DOWNTO 0);
     L551              :in std_logic_vector(8 DOWNTO 0);
     L552              :in std_logic_vector(8 DOWNTO 0);
     L553              :in std_logic_vector(8 DOWNTO 0);
     L554              :in std_logic_vector(8 DOWNTO 0);
     L555              :in std_logic_vector(8 DOWNTO 0);
     L556              :in std_logic_vector(8 DOWNTO 0);
     L557              :in std_logic_vector(8 DOWNTO 0);
     L558              :in std_logic_vector(8 DOWNTO 0);
     L559              :in std_logic_vector(8 DOWNTO 0);
     L560              :in std_logic_vector(8 DOWNTO 0);
     L561              :in std_logic_vector(8 DOWNTO 0);
     L562              :in std_logic_vector(8 DOWNTO 0);
     L563              :in std_logic_vector(8 DOWNTO 0);
     L564              :in std_logic_vector(8 DOWNTO 0);
     L565              :in std_logic_vector(8 DOWNTO 0);
     L566              :in std_logic_vector(8 DOWNTO 0);
     L567              :in std_logic_vector(8 DOWNTO 0);
     L568              :in std_logic_vector(8 DOWNTO 0);
     L569              :in std_logic_vector(8 DOWNTO 0);
     L570              :in std_logic_vector(8 DOWNTO 0);
     L571              :in std_logic_vector(8 DOWNTO 0);
     L572              :in std_logic_vector(8 DOWNTO 0);
     L573              :in std_logic_vector(8 DOWNTO 0);
     L574              :in std_logic_vector(8 DOWNTO 0);
     L575              :in std_logic_vector(8 DOWNTO 0);
     L576              :in std_logic_vector(8 DOWNTO 0);
     L577              :in std_logic_vector(8 DOWNTO 0);
     L578              :in std_logic_vector(8 DOWNTO 0);
     L579              :in std_logic_vector(8 DOWNTO 0);
     L580              :in std_logic_vector(8 DOWNTO 0);
     L581              :in std_logic_vector(8 DOWNTO 0);
     L582              :in std_logic_vector(8 DOWNTO 0);
     L583              :in std_logic_vector(8 DOWNTO 0);
     L584              :in std_logic_vector(8 DOWNTO 0);
     L585              :in std_logic_vector(8 DOWNTO 0);
     L586              :in std_logic_vector(8 DOWNTO 0);
     L587              :in std_logic_vector(8 DOWNTO 0);
     L588              :in std_logic_vector(8 DOWNTO 0);
     L589              :in std_logic_vector(8 DOWNTO 0);
     L590              :in std_logic_vector(8 DOWNTO 0);
     L591              :in std_logic_vector(8 DOWNTO 0);
     L592              :in std_logic_vector(8 DOWNTO 0);
     L593              :in std_logic_vector(8 DOWNTO 0);
     L594              :in std_logic_vector(8 DOWNTO 0);
     L595              :in std_logic_vector(8 DOWNTO 0);
     L596              :in std_logic_vector(8 DOWNTO 0);
     L597              :in std_logic_vector(8 DOWNTO 0);
     L598              :in std_logic_vector(8 DOWNTO 0);
     L599              :in std_logic_vector(8 DOWNTO 0);
     L600              :in std_logic_vector(8 DOWNTO 0);
     L601              :in std_logic_vector(8 DOWNTO 0);
     L602              :in std_logic_vector(8 DOWNTO 0);
     L603              :in std_logic_vector(8 DOWNTO 0);
     L604              :in std_logic_vector(8 DOWNTO 0);
     L605              :in std_logic_vector(8 DOWNTO 0);
     L606              :in std_logic_vector(8 DOWNTO 0);
     L607              :in std_logic_vector(8 DOWNTO 0);
     L608              :in std_logic_vector(8 DOWNTO 0);
     L609              :in std_logic_vector(8 DOWNTO 0);
     L610              :in std_logic_vector(8 DOWNTO 0);
     L611              :in std_logic_vector(8 DOWNTO 0);
     L612              :in std_logic_vector(8 DOWNTO 0);
     L613              :in std_logic_vector(8 DOWNTO 0);
     L614              :in std_logic_vector(8 DOWNTO 0);
     L615              :in std_logic_vector(8 DOWNTO 0);
     L616              :in std_logic_vector(8 DOWNTO 0);
     L617              :in std_logic_vector(8 DOWNTO 0);
     L618              :in std_logic_vector(8 DOWNTO 0);
     L619              :in std_logic_vector(8 DOWNTO 0);
     L620              :in std_logic_vector(8 DOWNTO 0);
     L621              :in std_logic_vector(8 DOWNTO 0);
     L622              :in std_logic_vector(8 DOWNTO 0);
     L623              :in std_logic_vector(8 DOWNTO 0);
     L624              :in std_logic_vector(8 DOWNTO 0);
     L625              :in std_logic_vector(8 DOWNTO 0);
     L626              :in std_logic_vector(8 DOWNTO 0);
     L627              :in std_logic_vector(8 DOWNTO 0);
     L628              :in std_logic_vector(8 DOWNTO 0);
     L629              :in std_logic_vector(8 DOWNTO 0);
     L630              :in std_logic_vector(8 DOWNTO 0);
     L631              :in std_logic_vector(8 DOWNTO 0);
     L632              :in std_logic_vector(8 DOWNTO 0);
     L633              :in std_logic_vector(8 DOWNTO 0);
     L634              :in std_logic_vector(8 DOWNTO 0);
     L635              :in std_logic_vector(8 DOWNTO 0);
     L636              :in std_logic_vector(8 DOWNTO 0);
     L637              :in std_logic_vector(8 DOWNTO 0);
     L638              :in std_logic_vector(8 DOWNTO 0);
     L639              :in std_logic_vector(8 DOWNTO 0);
     L640              :in std_logic_vector(8 DOWNTO 0);
     L641              :in std_logic_vector(8 DOWNTO 0);
     L642              :in std_logic_vector(8 DOWNTO 0);
     L643              :in std_logic_vector(8 DOWNTO 0);
     L644              :in std_logic_vector(8 DOWNTO 0);
     L645              :in std_logic_vector(8 DOWNTO 0);
     L646              :in std_logic_vector(8 DOWNTO 0);
     L647              :in std_logic_vector(8 DOWNTO 0);
     L648              :in std_logic_vector(8 DOWNTO 0);
     L649              :in std_logic_vector(8 DOWNTO 0);
     L650              :in std_logic_vector(8 DOWNTO 0);
     L651              :in std_logic_vector(8 DOWNTO 0);
     L652              :in std_logic_vector(8 DOWNTO 0);
     L653              :in std_logic_vector(8 DOWNTO 0);
     L654              :in std_logic_vector(8 DOWNTO 0);
     L655              :in std_logic_vector(8 DOWNTO 0);
     L656              :in std_logic_vector(8 DOWNTO 0);
     L657              :in std_logic_vector(8 DOWNTO 0);
     L658              :in std_logic_vector(8 DOWNTO 0);
     L659              :in std_logic_vector(8 DOWNTO 0);
     L660              :in std_logic_vector(8 DOWNTO 0);
     L661              :in std_logic_vector(8 DOWNTO 0);
     L662              :in std_logic_vector(8 DOWNTO 0);
     L663              :in std_logic_vector(8 DOWNTO 0);
     L664              :in std_logic_vector(8 DOWNTO 0);
     L665              :in std_logic_vector(8 DOWNTO 0);
     L666              :in std_logic_vector(8 DOWNTO 0);
     L667              :in std_logic_vector(8 DOWNTO 0);
     L668              :in std_logic_vector(8 DOWNTO 0);
     L669              :in std_logic_vector(8 DOWNTO 0);
     L670              :in std_logic_vector(8 DOWNTO 0);
     L671              :in std_logic_vector(8 DOWNTO 0);
     L672              :in std_logic_vector(8 DOWNTO 0);
     L673              :in std_logic_vector(8 DOWNTO 0);
     L674              :in std_logic_vector(8 DOWNTO 0);
     L675              :in std_logic_vector(8 DOWNTO 0);
     L676              :in std_logic_vector(8 DOWNTO 0);
     L677              :in std_logic_vector(8 DOWNTO 0);
     L678              :in std_logic_vector(8 DOWNTO 0);
     L679              :in std_logic_vector(8 DOWNTO 0);
     L680              :in std_logic_vector(8 DOWNTO 0);
     L681              :in std_logic_vector(8 DOWNTO 0);
     L682              :in std_logic_vector(8 DOWNTO 0);
     L683              :in std_logic_vector(8 DOWNTO 0);
     L684              :in std_logic_vector(8 DOWNTO 0);
     L685              :in std_logic_vector(8 DOWNTO 0);
     L686              :in std_logic_vector(8 DOWNTO 0);
     L687              :in std_logic_vector(8 DOWNTO 0);
     L688              :in std_logic_vector(8 DOWNTO 0);
     L689              :in std_logic_vector(8 DOWNTO 0);
     L690              :in std_logic_vector(8 DOWNTO 0);
     L691              :in std_logic_vector(8 DOWNTO 0);
     L692              :in std_logic_vector(8 DOWNTO 0);
     L693              :in std_logic_vector(8 DOWNTO 0);
     L694              :in std_logic_vector(8 DOWNTO 0);
     L695              :in std_logic_vector(8 DOWNTO 0);
     L696              :in std_logic_vector(8 DOWNTO 0);
     L697              :in std_logic_vector(8 DOWNTO 0);
     L698              :in std_logic_vector(8 DOWNTO 0);
     L699              :in std_logic_vector(8 DOWNTO 0);
     L700              :in std_logic_vector(8 DOWNTO 0);
     L701              :in std_logic_vector(8 DOWNTO 0);
     L702              :in std_logic_vector(8 DOWNTO 0);
     L703              :in std_logic_vector(8 DOWNTO 0);
     L704              :in std_logic_vector(8 DOWNTO 0);
     L705              :in std_logic_vector(8 DOWNTO 0);
     L706              :in std_logic_vector(8 DOWNTO 0);
     L707              :in std_logic_vector(8 DOWNTO 0);
     L708              :in std_logic_vector(8 DOWNTO 0);
     L709              :in std_logic_vector(8 DOWNTO 0);
     L710              :in std_logic_vector(8 DOWNTO 0);
     L711              :in std_logic_vector(8 DOWNTO 0);
     L712              :in std_logic_vector(8 DOWNTO 0);
     L713              :in std_logic_vector(8 DOWNTO 0);
     L714              :in std_logic_vector(8 DOWNTO 0);
     L715              :in std_logic_vector(8 DOWNTO 0);
     L716              :in std_logic_vector(8 DOWNTO 0);
     L717              :in std_logic_vector(8 DOWNTO 0);
     L718              :in std_logic_vector(8 DOWNTO 0);
     L719              :in std_logic_vector(8 DOWNTO 0);
     L720              :in std_logic_vector(8 DOWNTO 0);
     L721              :in std_logic_vector(8 DOWNTO 0);
     L722              :in std_logic_vector(8 DOWNTO 0);
     L723              :in std_logic_vector(8 DOWNTO 0);
     L724              :in std_logic_vector(8 DOWNTO 0);
     L725              :in std_logic_vector(8 DOWNTO 0);
     L726              :in std_logic_vector(8 DOWNTO 0);
     L727              :in std_logic_vector(8 DOWNTO 0);
     L728              :in std_logic_vector(8 DOWNTO 0);
     L729              :in std_logic_vector(8 DOWNTO 0);
     L730              :in std_logic_vector(8 DOWNTO 0);
     L731              :in std_logic_vector(8 DOWNTO 0);
     L732              :in std_logic_vector(8 DOWNTO 0);
     L733              :in std_logic_vector(8 DOWNTO 0);
     L734              :in std_logic_vector(8 DOWNTO 0);
     L735              :in std_logic_vector(8 DOWNTO 0);
     L736              :in std_logic_vector(8 DOWNTO 0);
     L737              :in std_logic_vector(8 DOWNTO 0);
     L738              :in std_logic_vector(8 DOWNTO 0);
     L739              :in std_logic_vector(8 DOWNTO 0);
     L740              :in std_logic_vector(8 DOWNTO 0);
     L741              :in std_logic_vector(8 DOWNTO 0);
     L742              :in std_logic_vector(8 DOWNTO 0);
     L743              :in std_logic_vector(8 DOWNTO 0);
     L744              :in std_logic_vector(8 DOWNTO 0);
     L745              :in std_logic_vector(8 DOWNTO 0);
     L746              :in std_logic_vector(8 DOWNTO 0);
     L747              :in std_logic_vector(8 DOWNTO 0);
     L748              :in std_logic_vector(8 DOWNTO 0);
     L749              :in std_logic_vector(8 DOWNTO 0);
     L750              :in std_logic_vector(8 DOWNTO 0);
     L751              :in std_logic_vector(8 DOWNTO 0);
     L752              :in std_logic_vector(8 DOWNTO 0);
     L753              :in std_logic_vector(8 DOWNTO 0);
     L754              :in std_logic_vector(8 DOWNTO 0);
     L755              :in std_logic_vector(8 DOWNTO 0);
     L756              :in std_logic_vector(8 DOWNTO 0);
     L757              :in std_logic_vector(8 DOWNTO 0);
     L758              :in std_logic_vector(8 DOWNTO 0);
     L759              :in std_logic_vector(8 DOWNTO 0);
     L760              :in std_logic_vector(8 DOWNTO 0);
     L761              :in std_logic_vector(8 DOWNTO 0);
     L762              :in std_logic_vector(8 DOWNTO 0);
     L763              :in std_logic_vector(8 DOWNTO 0);
     L764              :in std_logic_vector(8 DOWNTO 0);
     L765              :in std_logic_vector(8 DOWNTO 0);
     L766              :in std_logic_vector(8 DOWNTO 0);
     L767              :in std_logic_vector(8 DOWNTO 0);
     L768              :in std_logic_vector(8 DOWNTO 0);
     L769              :in std_logic_vector(8 DOWNTO 0);
     L770              :in std_logic_vector(8 DOWNTO 0);
     L771              :in std_logic_vector(8 DOWNTO 0);
     L772              :in std_logic_vector(8 DOWNTO 0);
     L773              :in std_logic_vector(8 DOWNTO 0);
     L774              :in std_logic_vector(8 DOWNTO 0);
     L775              :in std_logic_vector(8 DOWNTO 0);
     L776              :in std_logic_vector(8 DOWNTO 0);
     L777              :in std_logic_vector(8 DOWNTO 0);
     L778              :in std_logic_vector(8 DOWNTO 0);
     L779              :in std_logic_vector(8 DOWNTO 0);
     L780              :in std_logic_vector(8 DOWNTO 0);
     L781              :in std_logic_vector(8 DOWNTO 0);
     L782              :in std_logic_vector(8 DOWNTO 0);
     L783              :in std_logic_vector(8 DOWNTO 0);
     L784              :in std_logic_vector(8 DOWNTO 0);
     L785              :in std_logic_vector(8 DOWNTO 0);
     L786              :in std_logic_vector(8 DOWNTO 0);
     L787              :in std_logic_vector(8 DOWNTO 0);
     L788              :in std_logic_vector(8 DOWNTO 0);
     L789              :in std_logic_vector(8 DOWNTO 0);
     L790              :in std_logic_vector(8 DOWNTO 0);
     L791              :in std_logic_vector(8 DOWNTO 0);
     L792              :in std_logic_vector(8 DOWNTO 0);
     L793              :in std_logic_vector(8 DOWNTO 0);
     L794              :in std_logic_vector(8 DOWNTO 0);
     L795              :in std_logic_vector(8 DOWNTO 0);
     L796              :in std_logic_vector(8 DOWNTO 0);
     L797              :in std_logic_vector(8 DOWNTO 0);
     L798              :in std_logic_vector(8 DOWNTO 0);
     L799              :in std_logic_vector(8 DOWNTO 0);
     L800              :in std_logic_vector(8 DOWNTO 0);
     L801              :in std_logic_vector(8 DOWNTO 0);
     L802              :in std_logic_vector(8 DOWNTO 0);
     L803              :in std_logic_vector(8 DOWNTO 0);
     L804              :in std_logic_vector(8 DOWNTO 0);
     L805              :in std_logic_vector(8 DOWNTO 0);
     L806              :in std_logic_vector(8 DOWNTO 0);
     L807              :in std_logic_vector(8 DOWNTO 0);
     L808              :in std_logic_vector(8 DOWNTO 0);
     L809              :in std_logic_vector(8 DOWNTO 0);
     L810              :in std_logic_vector(8 DOWNTO 0);
     L811              :in std_logic_vector(8 DOWNTO 0);
     L812              :in std_logic_vector(8 DOWNTO 0);
     L813              :in std_logic_vector(8 DOWNTO 0);
     L814              :in std_logic_vector(8 DOWNTO 0);
     L815              :in std_logic_vector(8 DOWNTO 0);
     L816              :in std_logic_vector(8 DOWNTO 0);
     L817              :in std_logic_vector(8 DOWNTO 0);
     L818              :in std_logic_vector(8 DOWNTO 0);
     L819              :in std_logic_vector(8 DOWNTO 0);
     L820              :in std_logic_vector(8 DOWNTO 0);
     L821              :in std_logic_vector(8 DOWNTO 0);
     L822              :in std_logic_vector(8 DOWNTO 0);
     L823              :in std_logic_vector(8 DOWNTO 0);
     L824              :in std_logic_vector(8 DOWNTO 0);
     L825              :in std_logic_vector(8 DOWNTO 0);
     L826              :in std_logic_vector(8 DOWNTO 0);
     L827              :in std_logic_vector(8 DOWNTO 0);
     L828              :in std_logic_vector(8 DOWNTO 0);
     L829              :in std_logic_vector(8 DOWNTO 0);
     L830              :in std_logic_vector(8 DOWNTO 0);
     L831              :in std_logic_vector(8 DOWNTO 0);
     L832              :in std_logic_vector(8 DOWNTO 0);
     L833              :in std_logic_vector(8 DOWNTO 0);
     L834              :in std_logic_vector(8 DOWNTO 0);
     L835              :in std_logic_vector(8 DOWNTO 0);
     L836              :in std_logic_vector(8 DOWNTO 0);
     L837              :in std_logic_vector(8 DOWNTO 0);
     L838              :in std_logic_vector(8 DOWNTO 0);
     L839              :in std_logic_vector(8 DOWNTO 0);
     L840              :in std_logic_vector(8 DOWNTO 0);
     L841              :in std_logic_vector(8 DOWNTO 0);
     L842              :in std_logic_vector(8 DOWNTO 0);
     L843              :in std_logic_vector(8 DOWNTO 0);
     L844              :in std_logic_vector(8 DOWNTO 0);
     L845              :in std_logic_vector(8 DOWNTO 0);
     L846              :in std_logic_vector(8 DOWNTO 0);
     L847              :in std_logic_vector(8 DOWNTO 0);
     L848              :in std_logic_vector(8 DOWNTO 0);
     L849              :in std_logic_vector(8 DOWNTO 0);
     L850              :in std_logic_vector(8 DOWNTO 0);
     L851              :in std_logic_vector(8 DOWNTO 0);
     L852              :in std_logic_vector(8 DOWNTO 0);
     L853              :in std_logic_vector(8 DOWNTO 0);
     L854              :in std_logic_vector(8 DOWNTO 0);
     L855              :in std_logic_vector(8 DOWNTO 0);
     L856              :in std_logic_vector(8 DOWNTO 0);
     L857              :in std_logic_vector(8 DOWNTO 0);
     L858              :in std_logic_vector(8 DOWNTO 0);
     L859              :in std_logic_vector(8 DOWNTO 0);
     L860              :in std_logic_vector(8 DOWNTO 0);
     L861              :in std_logic_vector(8 DOWNTO 0);
     L862              :in std_logic_vector(8 DOWNTO 0);
     L863              :in std_logic_vector(8 DOWNTO 0);
     L864              :in std_logic_vector(8 DOWNTO 0);
     L865              :in std_logic_vector(8 DOWNTO 0);
     L866              :in std_logic_vector(8 DOWNTO 0);
     L867              :in std_logic_vector(8 DOWNTO 0);
     L868              :in std_logic_vector(8 DOWNTO 0);
     L869              :in std_logic_vector(8 DOWNTO 0);
     L870              :in std_logic_vector(8 DOWNTO 0);
     L871              :in std_logic_vector(8 DOWNTO 0);
     L872              :in std_logic_vector(8 DOWNTO 0);
     L873              :in std_logic_vector(8 DOWNTO 0);
     L874              :in std_logic_vector(8 DOWNTO 0);
     L875              :in std_logic_vector(8 DOWNTO 0);
     L876              :in std_logic_vector(8 DOWNTO 0);
     L877              :in std_logic_vector(8 DOWNTO 0);
     L878              :in std_logic_vector(8 DOWNTO 0);
     L879              :in std_logic_vector(8 DOWNTO 0);
     L880              :in std_logic_vector(8 DOWNTO 0);
     L881              :in std_logic_vector(8 DOWNTO 0);
     L882              :in std_logic_vector(8 DOWNTO 0);
     L883              :in std_logic_vector(8 DOWNTO 0);
     L884              :in std_logic_vector(8 DOWNTO 0);
     L885              :in std_logic_vector(8 DOWNTO 0);
     L886              :in std_logic_vector(8 DOWNTO 0);
     L887              :in std_logic_vector(8 DOWNTO 0);
     L888              :in std_logic_vector(8 DOWNTO 0);
     L889              :in std_logic_vector(8 DOWNTO 0);
     L890              :in std_logic_vector(8 DOWNTO 0);
     L891              :in std_logic_vector(8 DOWNTO 0);
     L892              :in std_logic_vector(8 DOWNTO 0);
     L893              :in std_logic_vector(8 DOWNTO 0);
     L894              :in std_logic_vector(8 DOWNTO 0);
     L895              :in std_logic_vector(8 DOWNTO 0);
     L896              :in std_logic_vector(8 DOWNTO 0);
     L897              :in std_logic_vector(8 DOWNTO 0);
     L898              :in std_logic_vector(8 DOWNTO 0);
     L899              :in std_logic_vector(8 DOWNTO 0);
     L900              :in std_logic_vector(8 DOWNTO 0);
     L901              :in std_logic_vector(8 DOWNTO 0);
     L902              :in std_logic_vector(8 DOWNTO 0);
     L903              :in std_logic_vector(8 DOWNTO 0);
     L904              :in std_logic_vector(8 DOWNTO 0);
     L905              :in std_logic_vector(8 DOWNTO 0);
     L906              :in std_logic_vector(8 DOWNTO 0);
     L907              :in std_logic_vector(8 DOWNTO 0);
     L908              :in std_logic_vector(8 DOWNTO 0);
     L909              :in std_logic_vector(8 DOWNTO 0);
     L910              :in std_logic_vector(8 DOWNTO 0);
     L911              :in std_logic_vector(8 DOWNTO 0);
     L912              :in std_logic_vector(8 DOWNTO 0);
     L913              :in std_logic_vector(8 DOWNTO 0);
     L914              :in std_logic_vector(8 DOWNTO 0);
     L915              :in std_logic_vector(8 DOWNTO 0);
     L916              :in std_logic_vector(8 DOWNTO 0);
     L917              :in std_logic_vector(8 DOWNTO 0);
     L918              :in std_logic_vector(8 DOWNTO 0);
     L919              :in std_logic_vector(8 DOWNTO 0);
     L920              :in std_logic_vector(8 DOWNTO 0);
     L921              :in std_logic_vector(8 DOWNTO 0);
     L922              :in std_logic_vector(8 DOWNTO 0);
     L923              :in std_logic_vector(8 DOWNTO 0);
     L924              :in std_logic_vector(8 DOWNTO 0);
     L925              :in std_logic_vector(8 DOWNTO 0);
     L926              :in std_logic_vector(8 DOWNTO 0);
     L927              :in std_logic_vector(8 DOWNTO 0);
     L928              :in std_logic_vector(8 DOWNTO 0);
     L929              :in std_logic_vector(8 DOWNTO 0);
     L930              :in std_logic_vector(8 DOWNTO 0);
     L931              :in std_logic_vector(8 DOWNTO 0);
     L932              :in std_logic_vector(8 DOWNTO 0);
     L933              :in std_logic_vector(8 DOWNTO 0);
     L934              :in std_logic_vector(8 DOWNTO 0);
     L935              :in std_logic_vector(8 DOWNTO 0);
     L936              :in std_logic_vector(8 DOWNTO 0);
     L937              :in std_logic_vector(8 DOWNTO 0);
     L938              :in std_logic_vector(8 DOWNTO 0);
     L939              :in std_logic_vector(8 DOWNTO 0);
     L940              :in std_logic_vector(8 DOWNTO 0);
     L941              :in std_logic_vector(8 DOWNTO 0);
     L942              :in std_logic_vector(8 DOWNTO 0);
     L943              :in std_logic_vector(8 DOWNTO 0);
     L944              :in std_logic_vector(8 DOWNTO 0);
     L945              :in std_logic_vector(8 DOWNTO 0);
     L946              :in std_logic_vector(8 DOWNTO 0);
     L947              :in std_logic_vector(8 DOWNTO 0);
     L948              :in std_logic_vector(8 DOWNTO 0);
     L949              :in std_logic_vector(8 DOWNTO 0);
     L950              :in std_logic_vector(8 DOWNTO 0);
     L951              :in std_logic_vector(8 DOWNTO 0);
     L952              :in std_logic_vector(8 DOWNTO 0);
     L953              :in std_logic_vector(8 DOWNTO 0);
     L954              :in std_logic_vector(8 DOWNTO 0);
     L955              :in std_logic_vector(8 DOWNTO 0);
     L956              :in std_logic_vector(8 DOWNTO 0);
     L957              :in std_logic_vector(8 DOWNTO 0);
     L958              :in std_logic_vector(8 DOWNTO 0);
     L959              :in std_logic_vector(8 DOWNTO 0);
     L960              :in std_logic_vector(8 DOWNTO 0);
     L961              :in std_logic_vector(8 DOWNTO 0);
     L962              :in std_logic_vector(8 DOWNTO 0);
     L963              :in std_logic_vector(8 DOWNTO 0);
     L964              :in std_logic_vector(8 DOWNTO 0);
     L965              :in std_logic_vector(8 DOWNTO 0);
     L966              :in std_logic_vector(8 DOWNTO 0);
     L967              :in std_logic_vector(8 DOWNTO 0);
     L968              :in std_logic_vector(8 DOWNTO 0);
     L969              :in std_logic_vector(8 DOWNTO 0);
     L970              :in std_logic_vector(8 DOWNTO 0);
     L971              :in std_logic_vector(8 DOWNTO 0);
     L972              :in std_logic_vector(8 DOWNTO 0);
     L973              :in std_logic_vector(8 DOWNTO 0);
     L974              :in std_logic_vector(8 DOWNTO 0);
     L975              :in std_logic_vector(8 DOWNTO 0);
     L976              :in std_logic_vector(8 DOWNTO 0);
     L977              :in std_logic_vector(8 DOWNTO 0);
     L978              :in std_logic_vector(8 DOWNTO 0);
     L979              :in std_logic_vector(8 DOWNTO 0);
     L980              :in std_logic_vector(8 DOWNTO 0);
     L981              :in std_logic_vector(8 DOWNTO 0);
     L982              :in std_logic_vector(8 DOWNTO 0);
     L983              :in std_logic_vector(8 DOWNTO 0);
     L984              :in std_logic_vector(8 DOWNTO 0);
     L985              :in std_logic_vector(8 DOWNTO 0);
     L986              :in std_logic_vector(8 DOWNTO 0);
     L987              :in std_logic_vector(8 DOWNTO 0);
     L988              :in std_logic_vector(8 DOWNTO 0);
     L989              :in std_logic_vector(8 DOWNTO 0);
     L990              :in std_logic_vector(8 DOWNTO 0);
     L991              :in std_logic_vector(8 DOWNTO 0);
     L992              :in std_logic_vector(8 DOWNTO 0);
     L993              :in std_logic_vector(8 DOWNTO 0);
     L994              :in std_logic_vector(8 DOWNTO 0);
     L995              :in std_logic_vector(8 DOWNTO 0);
     L996              :in std_logic_vector(8 DOWNTO 0);
     L997              :in std_logic_vector(8 DOWNTO 0);
     L998              :in std_logic_vector(8 DOWNTO 0);
     L999              :in std_logic_vector(8 DOWNTO 0);
     L1000              :in std_logic_vector(8 DOWNTO 0);
     L1001              :in std_logic_vector(8 DOWNTO 0);
     L1002              :in std_logic_vector(8 DOWNTO 0);
     L1003              :in std_logic_vector(8 DOWNTO 0);
     L1004              :in std_logic_vector(8 DOWNTO 0);
     L1005              :in std_logic_vector(8 DOWNTO 0);
     L1006              :in std_logic_vector(8 DOWNTO 0);
     L1007              :in std_logic_vector(8 DOWNTO 0);
     L1008              :in std_logic_vector(8 DOWNTO 0);
     L1009              :in std_logic_vector(8 DOWNTO 0);
     L1010              :in std_logic_vector(8 DOWNTO 0);
     L1011              :in std_logic_vector(8 DOWNTO 0);
     L1012              :in std_logic_vector(8 DOWNTO 0);
     L1013              :in std_logic_vector(8 DOWNTO 0);
     L1014              :in std_logic_vector(8 DOWNTO 0);
     L1015              :in std_logic_vector(8 DOWNTO 0);
     L1016              :in std_logic_vector(8 DOWNTO 0);
     L1017              :in std_logic_vector(8 DOWNTO 0);
     L1018              :in std_logic_vector(8 DOWNTO 0);
     L1019              :in std_logic_vector(8 DOWNTO 0);
     L1020              :in std_logic_vector(8 DOWNTO 0);
     L1021              :in std_logic_vector(8 DOWNTO 0);
     L1022              :in std_logic_vector(8 DOWNTO 0);
     L1023              :in std_logic_vector(8 DOWNTO 0);
     L1024              :in std_logic_vector(8 DOWNTO 0);
     L1025              :in std_logic_vector(8 DOWNTO 0);
     L1026              :in std_logic_vector(8 DOWNTO 0);
     L1027              :in std_logic_vector(8 DOWNTO 0);
     L1028              :in std_logic_vector(8 DOWNTO 0);
     L1029              :in std_logic_vector(8 DOWNTO 0);
     L1030              :in std_logic_vector(8 DOWNTO 0);
     L1031              :in std_logic_vector(8 DOWNTO 0);
     L1032              :in std_logic_vector(8 DOWNTO 0);
     L1033              :in std_logic_vector(8 DOWNTO 0);
     L1034              :in std_logic_vector(8 DOWNTO 0);
     L1035              :in std_logic_vector(8 DOWNTO 0);
     L1036              :in std_logic_vector(8 DOWNTO 0);
     L1037              :in std_logic_vector(8 DOWNTO 0);
     L1038              :in std_logic_vector(8 DOWNTO 0);
     L1039              :in std_logic_vector(8 DOWNTO 0);
     L1040              :in std_logic_vector(8 DOWNTO 0);
     L1041              :in std_logic_vector(8 DOWNTO 0);
     L1042              :in std_logic_vector(8 DOWNTO 0);
     L1043              :in std_logic_vector(8 DOWNTO 0);
     L1044              :in std_logic_vector(8 DOWNTO 0);
     L1045              :in std_logic_vector(8 DOWNTO 0);
     L1046              :in std_logic_vector(8 DOWNTO 0);
     L1047              :in std_logic_vector(8 DOWNTO 0);
     L1048              :in std_logic_vector(8 DOWNTO 0);
     L1049              :in std_logic_vector(8 DOWNTO 0);
     L1050              :in std_logic_vector(8 DOWNTO 0);
     L1051              :in std_logic_vector(8 DOWNTO 0);
     L1052              :in std_logic_vector(8 DOWNTO 0);
     L1053              :in std_logic_vector(8 DOWNTO 0);
     L1054              :in std_logic_vector(8 DOWNTO 0);
     L1055              :in std_logic_vector(8 DOWNTO 0);
     L1056              :in std_logic_vector(8 DOWNTO 0);
     L1057              :in std_logic_vector(8 DOWNTO 0);
     L1058              :in std_logic_vector(8 DOWNTO 0);
     L1059              :in std_logic_vector(8 DOWNTO 0);
     L1060              :in std_logic_vector(8 DOWNTO 0);
     L1061              :in std_logic_vector(8 DOWNTO 0);
     L1062              :in std_logic_vector(8 DOWNTO 0);
     L1063              :in std_logic_vector(8 DOWNTO 0);
     L1064              :in std_logic_vector(8 DOWNTO 0);
     L1065              :in std_logic_vector(8 DOWNTO 0);
     L1066              :in std_logic_vector(8 DOWNTO 0);
     L1067              :in std_logic_vector(8 DOWNTO 0);
     L1068              :in std_logic_vector(8 DOWNTO 0);
     L1069              :in std_logic_vector(8 DOWNTO 0);
     L1070              :in std_logic_vector(8 DOWNTO 0);
     L1071              :in std_logic_vector(8 DOWNTO 0);
     L1072              :in std_logic_vector(8 DOWNTO 0);
     L1073              :in std_logic_vector(8 DOWNTO 0);
     L1074              :in std_logic_vector(8 DOWNTO 0);
     L1075              :in std_logic_vector(8 DOWNTO 0);
     L1076              :in std_logic_vector(8 DOWNTO 0);
     L1077              :in std_logic_vector(8 DOWNTO 0);
     L1078              :in std_logic_vector(8 DOWNTO 0);
     L1079              :in std_logic_vector(8 DOWNTO 0);
     L1080              :in std_logic_vector(8 DOWNTO 0);
     L1081              :in std_logic_vector(8 DOWNTO 0);
     L1082              :in std_logic_vector(8 DOWNTO 0);
     L1083              :in std_logic_vector(8 DOWNTO 0);
     L1084              :in std_logic_vector(8 DOWNTO 0);
     L1085              :in std_logic_vector(8 DOWNTO 0);
     L1086              :in std_logic_vector(8 DOWNTO 0);
     L1087              :in std_logic_vector(8 DOWNTO 0);
     L1088              :in std_logic_vector(8 DOWNTO 0);
     L1089              :in std_logic_vector(8 DOWNTO 0);
     L1090              :in std_logic_vector(8 DOWNTO 0);
     L1091              :in std_logic_vector(8 DOWNTO 0);
     L1092              :in std_logic_vector(8 DOWNTO 0);
     L1093              :in std_logic_vector(8 DOWNTO 0);
     L1094              :in std_logic_vector(8 DOWNTO 0);
     L1095              :in std_logic_vector(8 DOWNTO 0);
     L1096              :in std_logic_vector(8 DOWNTO 0);
     L1097              :in std_logic_vector(8 DOWNTO 0);
     L1098              :in std_logic_vector(8 DOWNTO 0);
     L1099              :in std_logic_vector(8 DOWNTO 0);
     L1100              :in std_logic_vector(8 DOWNTO 0);
     L1101              :in std_logic_vector(8 DOWNTO 0);
     L1102              :in std_logic_vector(8 DOWNTO 0);
     L1103              :in std_logic_vector(8 DOWNTO 0);
     L1104              :in std_logic_vector(8 DOWNTO 0);
     L1105              :in std_logic_vector(8 DOWNTO 0);
     L1106              :in std_logic_vector(8 DOWNTO 0);
     L1107              :in std_logic_vector(8 DOWNTO 0);
     L1108              :in std_logic_vector(8 DOWNTO 0);
     L1109              :in std_logic_vector(8 DOWNTO 0);
     L1110              :in std_logic_vector(8 DOWNTO 0);
     L1111              :in std_logic_vector(8 DOWNTO 0);
     L1112              :in std_logic_vector(8 DOWNTO 0);
     L1113              :in std_logic_vector(8 DOWNTO 0);
     L1114              :in std_logic_vector(8 DOWNTO 0);
     L1115              :in std_logic_vector(8 DOWNTO 0);
     L1116              :in std_logic_vector(8 DOWNTO 0);
     L1117              :in std_logic_vector(8 DOWNTO 0);
     L1118              :in std_logic_vector(8 DOWNTO 0);
     L1119              :in std_logic_vector(8 DOWNTO 0);
     L1120              :in std_logic_vector(8 DOWNTO 0);
     L1121              :in std_logic_vector(8 DOWNTO 0);
     L1122              :in std_logic_vector(8 DOWNTO 0);
     L1123              :in std_logic_vector(8 DOWNTO 0);
     L1124              :in std_logic_vector(8 DOWNTO 0);
     L1125              :in std_logic_vector(8 DOWNTO 0);
     L1126              :in std_logic_vector(8 DOWNTO 0);
     L1127              :in std_logic_vector(8 DOWNTO 0);
     L1128              :in std_logic_vector(8 DOWNTO 0);
     L1129              :in std_logic_vector(8 DOWNTO 0);
     L1130              :in std_logic_vector(8 DOWNTO 0);
     L1131              :in std_logic_vector(8 DOWNTO 0);
     L1132              :in std_logic_vector(8 DOWNTO 0);
     L1133              :in std_logic_vector(8 DOWNTO 0);
     L1134              :in std_logic_vector(8 DOWNTO 0);
     L1135              :in std_logic_vector(8 DOWNTO 0);
     L1136              :in std_logic_vector(8 DOWNTO 0);
     L1137              :in std_logic_vector(8 DOWNTO 0);
     L1138              :in std_logic_vector(8 DOWNTO 0);
     L1139              :in std_logic_vector(8 DOWNTO 0);
     L1140              :in std_logic_vector(8 DOWNTO 0);
     L1141              :in std_logic_vector(8 DOWNTO 0);
     L1142              :in std_logic_vector(8 DOWNTO 0);
     L1143              :in std_logic_vector(8 DOWNTO 0);
     L1144              :in std_logic_vector(8 DOWNTO 0);
     L1145              :in std_logic_vector(8 DOWNTO 0);
     L1146              :in std_logic_vector(8 DOWNTO 0);
     L1147              :in std_logic_vector(8 DOWNTO 0);
     L1148              :in std_logic_vector(8 DOWNTO 0);
     L1149              :in std_logic_vector(8 DOWNTO 0);
     L1150              :in std_logic_vector(8 DOWNTO 0);
     L1151              :in std_logic_vector(8 DOWNTO 0);
     L1152              :in std_logic_vector(8 DOWNTO 0);
     L1153              :in std_logic_vector(8 DOWNTO 0);
     L1154              :in std_logic_vector(8 DOWNTO 0);
     L1155              :in std_logic_vector(8 DOWNTO 0);
     L1156              :in std_logic_vector(8 DOWNTO 0);
     L1157              :in std_logic_vector(8 DOWNTO 0);
     L1158              :in std_logic_vector(8 DOWNTO 0);
     L1159              :in std_logic_vector(8 DOWNTO 0);
     L1160              :in std_logic_vector(8 DOWNTO 0);
     L1161              :in std_logic_vector(8 DOWNTO 0);
     L1162              :in std_logic_vector(8 DOWNTO 0);
     L1163              :in std_logic_vector(8 DOWNTO 0);
     L1164              :in std_logic_vector(8 DOWNTO 0);
     L1165              :in std_logic_vector(8 DOWNTO 0);
     L1166              :in std_logic_vector(8 DOWNTO 0);
     L1167              :in std_logic_vector(8 DOWNTO 0);
     L1168              :in std_logic_vector(8 DOWNTO 0);
     L1169              :in std_logic_vector(8 DOWNTO 0);
     L1170              :in std_logic_vector(8 DOWNTO 0);
     L1171              :in std_logic_vector(8 DOWNTO 0);
     L1172              :in std_logic_vector(8 DOWNTO 0);
     L1173              :in std_logic_vector(8 DOWNTO 0);
     L1174              :in std_logic_vector(8 DOWNTO 0);
     L1175              :in std_logic_vector(8 DOWNTO 0);
     L1176              :in std_logic_vector(8 DOWNTO 0);
     L1177              :in std_logic_vector(8 DOWNTO 0);
     L1178              :in std_logic_vector(8 DOWNTO 0);
     L1179              :in std_logic_vector(8 DOWNTO 0);
     L1180              :in std_logic_vector(8 DOWNTO 0);
     L1181              :in std_logic_vector(8 DOWNTO 0);
     L1182              :in std_logic_vector(8 DOWNTO 0);
     L1183              :in std_logic_vector(8 DOWNTO 0);
     L1184              :in std_logic_vector(8 DOWNTO 0);
     L1185              :in std_logic_vector(8 DOWNTO 0);
     L1186              :in std_logic_vector(8 DOWNTO 0);
     L1187              :in std_logic_vector(8 DOWNTO 0);
     L1188              :in std_logic_vector(8 DOWNTO 0);
     L1189              :in std_logic_vector(8 DOWNTO 0);
     L1190              :in std_logic_vector(8 DOWNTO 0);
     L1191              :in std_logic_vector(8 DOWNTO 0);
     L1192              :in std_logic_vector(8 DOWNTO 0);
     L1193              :in std_logic_vector(8 DOWNTO 0);
     L1194              :in std_logic_vector(8 DOWNTO 0);
     L1195              :in std_logic_vector(8 DOWNTO 0);
     L1196              :in std_logic_vector(8 DOWNTO 0);
     L1197              :in std_logic_vector(8 DOWNTO 0);
     L1198              :in std_logic_vector(8 DOWNTO 0);
     L1199              :in std_logic_vector(8 DOWNTO 0);
     L1200              :in std_logic_vector(8 DOWNTO 0);
     L1201              :in std_logic_vector(8 DOWNTO 0);
     L1202              :in std_logic_vector(8 DOWNTO 0);
     L1203              :in std_logic_vector(8 DOWNTO 0);
     L1204              :in std_logic_vector(8 DOWNTO 0);
     L1205              :in std_logic_vector(8 DOWNTO 0);
     L1206              :in std_logic_vector(8 DOWNTO 0);
     L1207              :in std_logic_vector(8 DOWNTO 0);
     L1208              :in std_logic_vector(8 DOWNTO 0);
     L1209              :in std_logic_vector(8 DOWNTO 0);
     L1210              :in std_logic_vector(8 DOWNTO 0);
     L1211              :in std_logic_vector(8 DOWNTO 0);
     L1212              :in std_logic_vector(8 DOWNTO 0);
     L1213              :in std_logic_vector(8 DOWNTO 0);
     L1214              :in std_logic_vector(8 DOWNTO 0);
     L1215              :in std_logic_vector(8 DOWNTO 0);
     L1216              :in std_logic_vector(8 DOWNTO 0);
     L1217              :in std_logic_vector(8 DOWNTO 0);
     L1218              :in std_logic_vector(8 DOWNTO 0);
     L1219              :in std_logic_vector(8 DOWNTO 0);
     L1220              :in std_logic_vector(8 DOWNTO 0);
     L1221              :in std_logic_vector(8 DOWNTO 0);
     L1222              :in std_logic_vector(8 DOWNTO 0);
     L1223              :in std_logic_vector(8 DOWNTO 0);
     L1224              :in std_logic_vector(8 DOWNTO 0);
     L1225              :in std_logic_vector(8 DOWNTO 0);
     L1226              :in std_logic_vector(8 DOWNTO 0);
     L1227              :in std_logic_vector(8 DOWNTO 0);
     L1228              :in std_logic_vector(8 DOWNTO 0);
     L1229              :in std_logic_vector(8 DOWNTO 0);
     L1230              :in std_logic_vector(8 DOWNTO 0);
     L1231              :in std_logic_vector(8 DOWNTO 0);
     L1232              :in std_logic_vector(8 DOWNTO 0);
     L1233              :in std_logic_vector(8 DOWNTO 0);
     L1234              :in std_logic_vector(8 DOWNTO 0);
     L1235              :in std_logic_vector(8 DOWNTO 0);
     L1236              :in std_logic_vector(8 DOWNTO 0);
     L1237              :in std_logic_vector(8 DOWNTO 0);
     L1238              :in std_logic_vector(8 DOWNTO 0);
     L1239              :in std_logic_vector(8 DOWNTO 0);
     L1240              :in std_logic_vector(8 DOWNTO 0);
     L1241              :in std_logic_vector(8 DOWNTO 0);
     L1242              :in std_logic_vector(8 DOWNTO 0);
     L1243              :in std_logic_vector(8 DOWNTO 0);
     L1244              :in std_logic_vector(8 DOWNTO 0);
     L1245              :in std_logic_vector(8 DOWNTO 0);
     L1246              :in std_logic_vector(8 DOWNTO 0);
     L1247              :in std_logic_vector(8 DOWNTO 0);
     L1248              :in std_logic_vector(8 DOWNTO 0);
     L1249              :in std_logic_vector(8 DOWNTO 0);
     L1250              :in std_logic_vector(8 DOWNTO 0);
     L1251              :in std_logic_vector(8 DOWNTO 0);
     L1252              :in std_logic_vector(8 DOWNTO 0);
     L1253              :in std_logic_vector(8 DOWNTO 0);
     L1254              :in std_logic_vector(8 DOWNTO 0);
     L1255              :in std_logic_vector(8 DOWNTO 0);
     L1256              :in std_logic_vector(8 DOWNTO 0);
     L1257              :in std_logic_vector(8 DOWNTO 0);
     L1258              :in std_logic_vector(8 DOWNTO 0);
     L1259              :in std_logic_vector(8 DOWNTO 0);
     L1260              :in std_logic_vector(8 DOWNTO 0);
     L1261              :in std_logic_vector(8 DOWNTO 0);
     L1262              :in std_logic_vector(8 DOWNTO 0);
     L1263              :in std_logic_vector(8 DOWNTO 0);
     L1264              :in std_logic_vector(8 DOWNTO 0);
     L1265              :in std_logic_vector(8 DOWNTO 0);
     L1266              :in std_logic_vector(8 DOWNTO 0);
     L1267              :in std_logic_vector(8 DOWNTO 0);
     L1268              :in std_logic_vector(8 DOWNTO 0);
     L1269              :in std_logic_vector(8 DOWNTO 0);
     L1270              :in std_logic_vector(8 DOWNTO 0);
     L1271              :in std_logic_vector(8 DOWNTO 0);
     L1272              :in std_logic_vector(8 DOWNTO 0);
     L1273              :in std_logic_vector(8 DOWNTO 0);
     L1274              :in std_logic_vector(8 DOWNTO 0);
     L1275              :in std_logic_vector(8 DOWNTO 0);
     L1276              :in std_logic_vector(8 DOWNTO 0);
     L1277              :in std_logic_vector(8 DOWNTO 0);
     L1278              :in std_logic_vector(8 DOWNTO 0);
     L1279              :in std_logic_vector(8 DOWNTO 0);
     L1280              :in std_logic_vector(8 DOWNTO 0);
     L1281              :in std_logic_vector(8 DOWNTO 0);
     L1282              :in std_logic_vector(8 DOWNTO 0);
     L1283              :in std_logic_vector(8 DOWNTO 0);
     L1284              :in std_logic_vector(8 DOWNTO 0);
     L1285              :in std_logic_vector(8 DOWNTO 0);
     L1286              :in std_logic_vector(8 DOWNTO 0);
     L1287              :in std_logic_vector(8 DOWNTO 0);
     L1288              :in std_logic_vector(8 DOWNTO 0);
     L1289              :in std_logic_vector(8 DOWNTO 0);
     L1290              :in std_logic_vector(8 DOWNTO 0);
     L1291              :in std_logic_vector(8 DOWNTO 0);
     L1292              :in std_logic_vector(8 DOWNTO 0);
     L1293              :in std_logic_vector(8 DOWNTO 0);
     L1294              :in std_logic_vector(8 DOWNTO 0);
     L1295              :in std_logic_vector(8 DOWNTO 0);
     L1296              :in std_logic_vector(8 DOWNTO 0);
     L1297              :in std_logic_vector(8 DOWNTO 0);
     L1298              :in std_logic_vector(8 DOWNTO 0);
     L1299              :in std_logic_vector(8 DOWNTO 0);
     L1300              :in std_logic_vector(8 DOWNTO 0);
     L1301              :in std_logic_vector(8 DOWNTO 0);
     L1302              :in std_logic_vector(8 DOWNTO 0);
     L1303              :in std_logic_vector(8 DOWNTO 0);
     L1304              :in std_logic_vector(8 DOWNTO 0);
     L1305              :in std_logic_vector(8 DOWNTO 0);
     L1306              :in std_logic_vector(8 DOWNTO 0);
     L1307              :in std_logic_vector(8 DOWNTO 0);
     L1308              :in std_logic_vector(8 DOWNTO 0);
     L1309              :in std_logic_vector(8 DOWNTO 0);
     L1310              :in std_logic_vector(8 DOWNTO 0);
     L1311              :in std_logic_vector(8 DOWNTO 0);
     L1312              :in std_logic_vector(8 DOWNTO 0);
     L1313              :in std_logic_vector(8 DOWNTO 0);
     L1314              :in std_logic_vector(8 DOWNTO 0);
     L1315              :in std_logic_vector(8 DOWNTO 0);
     L1316              :in std_logic_vector(8 DOWNTO 0);
     L1317              :in std_logic_vector(8 DOWNTO 0);
     L1318              :in std_logic_vector(8 DOWNTO 0);
     L1319              :in std_logic_vector(8 DOWNTO 0);
     L1320              :in std_logic_vector(8 DOWNTO 0);
     L1321              :in std_logic_vector(8 DOWNTO 0);
     L1322              :in std_logic_vector(8 DOWNTO 0);
     L1323              :in std_logic_vector(8 DOWNTO 0);
     L1324              :in std_logic_vector(8 DOWNTO 0);
     L1325              :in std_logic_vector(8 DOWNTO 0);
     L1326              :in std_logic_vector(8 DOWNTO 0);
     L1327              :in std_logic_vector(8 DOWNTO 0);
     L1328              :in std_logic_vector(8 DOWNTO 0);
     L1329              :in std_logic_vector(8 DOWNTO 0);
     L1330              :in std_logic_vector(8 DOWNTO 0);
     L1331              :in std_logic_vector(8 DOWNTO 0);
     L1332              :in std_logic_vector(8 DOWNTO 0);
     L1333              :in std_logic_vector(8 DOWNTO 0);
     L1334              :in std_logic_vector(8 DOWNTO 0);
     L1335              :in std_logic_vector(8 DOWNTO 0);
     L1336              :in std_logic_vector(8 DOWNTO 0);
     L1337              :in std_logic_vector(8 DOWNTO 0);
     L1338              :in std_logic_vector(8 DOWNTO 0);
     L1339              :in std_logic_vector(8 DOWNTO 0);
     L1340              :in std_logic_vector(8 DOWNTO 0);
     L1341              :in std_logic_vector(8 DOWNTO 0);
     L1342              :in std_logic_vector(8 DOWNTO 0);
     L1343              :in std_logic_vector(8 DOWNTO 0);
     L1344              :in std_logic_vector(8 DOWNTO 0);
     L1345              :in std_logic_vector(8 DOWNTO 0);
     L1346              :in std_logic_vector(8 DOWNTO 0);
     L1347              :in std_logic_vector(8 DOWNTO 0);
     L1348              :in std_logic_vector(8 DOWNTO 0);
     L1349              :in std_logic_vector(8 DOWNTO 0);
     L1350              :in std_logic_vector(8 DOWNTO 0);
     L1351              :in std_logic_vector(8 DOWNTO 0);
     L1352              :in std_logic_vector(8 DOWNTO 0);
     L1353              :in std_logic_vector(8 DOWNTO 0);
     L1354              :in std_logic_vector(8 DOWNTO 0);
     L1355              :in std_logic_vector(8 DOWNTO 0);
     L1356              :in std_logic_vector(8 DOWNTO 0);
     L1357              :in std_logic_vector(8 DOWNTO 0);
     L1358              :in std_logic_vector(8 DOWNTO 0);
     L1359              :in std_logic_vector(8 DOWNTO 0);
     L1360              :in std_logic_vector(8 DOWNTO 0);
     L1361              :in std_logic_vector(8 DOWNTO 0);
     L1362              :in std_logic_vector(8 DOWNTO 0);
     L1363              :in std_logic_vector(8 DOWNTO 0);
     L1364              :in std_logic_vector(8 DOWNTO 0);
     L1365              :in std_logic_vector(8 DOWNTO 0);
     L1366              :in std_logic_vector(8 DOWNTO 0);
     L1367              :in std_logic_vector(8 DOWNTO 0);
     L1368              :in std_logic_vector(8 DOWNTO 0);
     L1369              :in std_logic_vector(8 DOWNTO 0);
     L1370              :in std_logic_vector(8 DOWNTO 0);
     L1371              :in std_logic_vector(8 DOWNTO 0);
     L1372              :in std_logic_vector(8 DOWNTO 0);
     L1373              :in std_logic_vector(8 DOWNTO 0);
     L1374              :in std_logic_vector(8 DOWNTO 0);
     L1375              :in std_logic_vector(8 DOWNTO 0);
     L1376              :in std_logic_vector(8 DOWNTO 0);
     L1377              :in std_logic_vector(8 DOWNTO 0);
     L1378              :in std_logic_vector(8 DOWNTO 0);
     L1379              :in std_logic_vector(8 DOWNTO 0);
     L1380              :in std_logic_vector(8 DOWNTO 0);
     L1381              :in std_logic_vector(8 DOWNTO 0);
     L1382              :in std_logic_vector(8 DOWNTO 0);
     L1383              :in std_logic_vector(8 DOWNTO 0);
     L1384              :in std_logic_vector(8 DOWNTO 0);
     L1385              :in std_logic_vector(8 DOWNTO 0);
     L1386              :in std_logic_vector(8 DOWNTO 0);
     L1387              :in std_logic_vector(8 DOWNTO 0);
     L1388              :in std_logic_vector(8 DOWNTO 0);
     L1389              :in std_logic_vector(8 DOWNTO 0);
     L1390              :in std_logic_vector(8 DOWNTO 0);
     L1391              :in std_logic_vector(8 DOWNTO 0);
     L1392              :in std_logic_vector(8 DOWNTO 0);
     L1393              :in std_logic_vector(8 DOWNTO 0);
     L1394              :in std_logic_vector(8 DOWNTO 0);
     L1395              :in std_logic_vector(8 DOWNTO 0);
     L1396              :in std_logic_vector(8 DOWNTO 0);
     L1397              :in std_logic_vector(8 DOWNTO 0);
     L1398              :in std_logic_vector(8 DOWNTO 0);
     L1399              :in std_logic_vector(8 DOWNTO 0);
     L1400              :in std_logic_vector(8 DOWNTO 0);
     L1401              :in std_logic_vector(8 DOWNTO 0);
     L1402              :in std_logic_vector(8 DOWNTO 0);
     L1403              :in std_logic_vector(8 DOWNTO 0);
     L1404              :in std_logic_vector(8 DOWNTO 0);
     L1405              :in std_logic_vector(8 DOWNTO 0);
     L1406              :in std_logic_vector(8 DOWNTO 0);
     L1407              :in std_logic_vector(8 DOWNTO 0);
     L1408              :in std_logic_vector(8 DOWNTO 0);
     L1409              :in std_logic_vector(8 DOWNTO 0);
     L1410              :in std_logic_vector(8 DOWNTO 0);
     L1411              :in std_logic_vector(8 DOWNTO 0);
     L1412              :in std_logic_vector(8 DOWNTO 0);
     L1413              :in std_logic_vector(8 DOWNTO 0);
     L1414              :in std_logic_vector(8 DOWNTO 0);
     L1415              :in std_logic_vector(8 DOWNTO 0);
     L1416              :in std_logic_vector(8 DOWNTO 0);
     L1417              :in std_logic_vector(8 DOWNTO 0);
     L1418              :in std_logic_vector(8 DOWNTO 0);
     L1419              :in std_logic_vector(8 DOWNTO 0);
     L1420              :in std_logic_vector(8 DOWNTO 0);
     L1421              :in std_logic_vector(8 DOWNTO 0);
     L1422              :in std_logic_vector(8 DOWNTO 0);
     L1423              :in std_logic_vector(8 DOWNTO 0);
     L1424              :in std_logic_vector(8 DOWNTO 0);
     L1425              :in std_logic_vector(8 DOWNTO 0);
     L1426              :in std_logic_vector(8 DOWNTO 0);
     L1427              :in std_logic_vector(8 DOWNTO 0);
     L1428              :in std_logic_vector(8 DOWNTO 0);
     L1429              :in std_logic_vector(8 DOWNTO 0);
     L1430              :in std_logic_vector(8 DOWNTO 0);
     L1431              :in std_logic_vector(8 DOWNTO 0);
     L1432              :in std_logic_vector(8 DOWNTO 0);
     L1433              :in std_logic_vector(8 DOWNTO 0);
     L1434              :in std_logic_vector(8 DOWNTO 0);
     L1435              :in std_logic_vector(8 DOWNTO 0);
     L1436              :in std_logic_vector(8 DOWNTO 0);
     L1437              :in std_logic_vector(8 DOWNTO 0);
     L1438              :in std_logic_vector(8 DOWNTO 0);
     L1439              :in std_logic_vector(8 DOWNTO 0);
     L1440              :in std_logic_vector(8 DOWNTO 0);
     L1441              :in std_logic_vector(8 DOWNTO 0);
     L1442              :in std_logic_vector(8 DOWNTO 0);
     L1443              :in std_logic_vector(8 DOWNTO 0);
     L1444              :in std_logic_vector(8 DOWNTO 0);
     L1445              :in std_logic_vector(8 DOWNTO 0);
     L1446              :in std_logic_vector(8 DOWNTO 0);
     L1447              :in std_logic_vector(8 DOWNTO 0);
     L1448              :in std_logic_vector(8 DOWNTO 0);
     L1449              :in std_logic_vector(8 DOWNTO 0);
     L1450              :in std_logic_vector(8 DOWNTO 0);
     L1451              :in std_logic_vector(8 DOWNTO 0);
     L1452              :in std_logic_vector(8 DOWNTO 0);
     L1453              :in std_logic_vector(8 DOWNTO 0);
     L1454              :in std_logic_vector(8 DOWNTO 0);
     L1455              :in std_logic_vector(8 DOWNTO 0);
     L1456              :in std_logic_vector(8 DOWNTO 0);
     L1457              :in std_logic_vector(8 DOWNTO 0);
     L1458              :in std_logic_vector(8 DOWNTO 0);
     L1459              :in std_logic_vector(8 DOWNTO 0);
     L1460              :in std_logic_vector(8 DOWNTO 0);
     L1461              :in std_logic_vector(8 DOWNTO 0);
     L1462              :in std_logic_vector(8 DOWNTO 0);
     L1463              :in std_logic_vector(8 DOWNTO 0);
     L1464              :in std_logic_vector(8 DOWNTO 0);
     L1465              :in std_logic_vector(8 DOWNTO 0);
     L1466              :in std_logic_vector(8 DOWNTO 0);
     L1467              :in std_logic_vector(8 DOWNTO 0);
     L1468              :in std_logic_vector(8 DOWNTO 0);
     L1469              :in std_logic_vector(8 DOWNTO 0);
     L1470              :in std_logic_vector(8 DOWNTO 0);
     L1471              :in std_logic_vector(8 DOWNTO 0);
     L1472              :in std_logic_vector(8 DOWNTO 0);
     L1473              :in std_logic_vector(8 DOWNTO 0);
     L1474              :in std_logic_vector(8 DOWNTO 0);
     L1475              :in std_logic_vector(8 DOWNTO 0);
     L1476              :in std_logic_vector(8 DOWNTO 0);
     L1477              :in std_logic_vector(8 DOWNTO 0);
     L1478              :in std_logic_vector(8 DOWNTO 0);
     L1479              :in std_logic_vector(8 DOWNTO 0);
     L1480              :in std_logic_vector(8 DOWNTO 0);
     L1481              :in std_logic_vector(8 DOWNTO 0);
     L1482              :in std_logic_vector(8 DOWNTO 0);
     L1483              :in std_logic_vector(8 DOWNTO 0);
     L1484              :in std_logic_vector(8 DOWNTO 0);
     L1485              :in std_logic_vector(8 DOWNTO 0);
     L1486              :in std_logic_vector(8 DOWNTO 0);
     L1487              :in std_logic_vector(8 DOWNTO 0);
     L1488              :in std_logic_vector(8 DOWNTO 0);
     L1489              :in std_logic_vector(8 DOWNTO 0);
     L1490              :in std_logic_vector(8 DOWNTO 0);
     L1491              :in std_logic_vector(8 DOWNTO 0);
     L1492              :in std_logic_vector(8 DOWNTO 0);
     L1493              :in std_logic_vector(8 DOWNTO 0);
     L1494              :in std_logic_vector(8 DOWNTO 0);
     L1495              :in std_logic_vector(8 DOWNTO 0);
     L1496              :in std_logic_vector(8 DOWNTO 0);
     L1497              :in std_logic_vector(8 DOWNTO 0);
     L1498              :in std_logic_vector(8 DOWNTO 0);
     L1499              :in std_logic_vector(8 DOWNTO 0);
     L1500              :in std_logic_vector(8 DOWNTO 0);
     L1501              :in std_logic_vector(8 DOWNTO 0);
     L1502              :in std_logic_vector(8 DOWNTO 0);
     L1503              :in std_logic_vector(8 DOWNTO 0);
     L1504              :in std_logic_vector(8 DOWNTO 0);
     L1505              :in std_logic_vector(8 DOWNTO 0);
     L1506              :in std_logic_vector(8 DOWNTO 0);
     L1507              :in std_logic_vector(8 DOWNTO 0);
     L1508              :in std_logic_vector(8 DOWNTO 0);
     L1509              :in std_logic_vector(8 DOWNTO 0);
     L1510              :in std_logic_vector(8 DOWNTO 0);
     L1511              :in std_logic_vector(8 DOWNTO 0);
     L1512              :in std_logic_vector(8 DOWNTO 0);
     L1513              :in std_logic_vector(8 DOWNTO 0);
     L1514              :in std_logic_vector(8 DOWNTO 0);
     L1515              :in std_logic_vector(8 DOWNTO 0);
     L1516              :in std_logic_vector(8 DOWNTO 0);
     L1517              :in std_logic_vector(8 DOWNTO 0);
     L1518              :in std_logic_vector(8 DOWNTO 0);
     L1519              :in std_logic_vector(8 DOWNTO 0);
     L1520              :in std_logic_vector(8 DOWNTO 0);
     L1521              :in std_logic_vector(8 DOWNTO 0);
     L1522              :in std_logic_vector(8 DOWNTO 0);
     L1523              :in std_logic_vector(8 DOWNTO 0);
     L1524              :in std_logic_vector(8 DOWNTO 0);
     L1525              :in std_logic_vector(8 DOWNTO 0);
     L1526              :in std_logic_vector(8 DOWNTO 0);
     L1527              :in std_logic_vector(8 DOWNTO 0);
     L1528              :in std_logic_vector(8 DOWNTO 0);
     L1529              :in std_logic_vector(8 DOWNTO 0);
     L1530              :in std_logic_vector(8 DOWNTO 0);
     L1531              :in std_logic_vector(8 DOWNTO 0);
     L1532              :in std_logic_vector(8 DOWNTO 0);
     L1533              :in std_logic_vector(8 DOWNTO 0);
     L1534              :in std_logic_vector(8 DOWNTO 0);
     L1535              :in std_logic_vector(8 DOWNTO 0);
     L1536              :in std_logic_vector(8 DOWNTO 0);
     L1537              :in std_logic_vector(8 DOWNTO 0);
     L1538              :in std_logic_vector(8 DOWNTO 0);
     L1539              :in std_logic_vector(8 DOWNTO 0);
     L1540              :in std_logic_vector(8 DOWNTO 0);
     L1541              :in std_logic_vector(8 DOWNTO 0);
     L1542              :in std_logic_vector(8 DOWNTO 0);
     L1543              :in std_logic_vector(8 DOWNTO 0);
     L1544              :in std_logic_vector(8 DOWNTO 0);
     L1545              :in std_logic_vector(8 DOWNTO 0);
     L1546              :in std_logic_vector(8 DOWNTO 0);
     L1547              :in std_logic_vector(8 DOWNTO 0);
     L1548              :in std_logic_vector(8 DOWNTO 0);
     L1549              :in std_logic_vector(8 DOWNTO 0);
     L1550              :in std_logic_vector(8 DOWNTO 0);
     L1551              :in std_logic_vector(8 DOWNTO 0);
     L1552              :in std_logic_vector(8 DOWNTO 0);
     L1553              :in std_logic_vector(8 DOWNTO 0);
     L1554              :in std_logic_vector(8 DOWNTO 0);
     L1555              :in std_logic_vector(8 DOWNTO 0);
     L1556              :in std_logic_vector(8 DOWNTO 0);
     L1557              :in std_logic_vector(8 DOWNTO 0);
     L1558              :in std_logic_vector(8 DOWNTO 0);
     L1559              :in std_logic_vector(8 DOWNTO 0);
     L1560              :in std_logic_vector(8 DOWNTO 0);
     L1561              :in std_logic_vector(8 DOWNTO 0);
     L1562              :in std_logic_vector(8 DOWNTO 0);
     L1563              :in std_logic_vector(8 DOWNTO 0);
     L1564              :in std_logic_vector(8 DOWNTO 0);
     L1565              :in std_logic_vector(8 DOWNTO 0);
     L1566              :in std_logic_vector(8 DOWNTO 0);
     L1567              :in std_logic_vector(8 DOWNTO 0);
     L1568              :in std_logic_vector(8 DOWNTO 0);
     L1569              :in std_logic_vector(8 DOWNTO 0);
     L1570              :in std_logic_vector(8 DOWNTO 0);
     L1571              :in std_logic_vector(8 DOWNTO 0);
     L1572              :in std_logic_vector(8 DOWNTO 0);
     L1573              :in std_logic_vector(8 DOWNTO 0);
     L1574              :in std_logic_vector(8 DOWNTO 0);
     L1575              :in std_logic_vector(8 DOWNTO 0);
     L1576              :in std_logic_vector(8 DOWNTO 0);
     L1577              :in std_logic_vector(8 DOWNTO 0);
     L1578              :in std_logic_vector(8 DOWNTO 0);
     L1579              :in std_logic_vector(8 DOWNTO 0);
     L1580              :in std_logic_vector(8 DOWNTO 0);
     L1581              :in std_logic_vector(8 DOWNTO 0);
     L1582              :in std_logic_vector(8 DOWNTO 0);
     L1583              :in std_logic_vector(8 DOWNTO 0);
     L1584              :in std_logic_vector(8 DOWNTO 0);
     L1585              :in std_logic_vector(8 DOWNTO 0);
     L1586              :in std_logic_vector(8 DOWNTO 0);
     L1587              :in std_logic_vector(8 DOWNTO 0);
     L1588              :in std_logic_vector(8 DOWNTO 0);
     L1589              :in std_logic_vector(8 DOWNTO 0);
     L1590              :in std_logic_vector(8 DOWNTO 0);
     L1591              :in std_logic_vector(8 DOWNTO 0);
     L1592              :in std_logic_vector(8 DOWNTO 0);
     L1593              :in std_logic_vector(8 DOWNTO 0);
     L1594              :in std_logic_vector(8 DOWNTO 0);
     L1595              :in std_logic_vector(8 DOWNTO 0);
     L1596              :in std_logic_vector(8 DOWNTO 0);
     L1597              :in std_logic_vector(8 DOWNTO 0);
     L1598              :in std_logic_vector(8 DOWNTO 0);
     L1599              :in std_logic_vector(8 DOWNTO 0);
     L1600              :in std_logic_vector(8 DOWNTO 0);
     L1601              :in std_logic_vector(8 DOWNTO 0);
     L1602              :in std_logic_vector(8 DOWNTO 0);
     L1603              :in std_logic_vector(8 DOWNTO 0);
     L1604              :in std_logic_vector(8 DOWNTO 0);
     L1605              :in std_logic_vector(8 DOWNTO 0);
     L1606              :in std_logic_vector(8 DOWNTO 0);
     L1607              :in std_logic_vector(8 DOWNTO 0);
     L1608              :in std_logic_vector(8 DOWNTO 0);
     L1609              :in std_logic_vector(8 DOWNTO 0);
     L1610              :in std_logic_vector(8 DOWNTO 0);
     L1611              :in std_logic_vector(8 DOWNTO 0);
     L1612              :in std_logic_vector(8 DOWNTO 0);
     L1613              :in std_logic_vector(8 DOWNTO 0);
     L1614              :in std_logic_vector(8 DOWNTO 0);
     L1615              :in std_logic_vector(8 DOWNTO 0);
     L1616              :in std_logic_vector(8 DOWNTO 0);
     L1617              :in std_logic_vector(8 DOWNTO 0);
     L1618              :in std_logic_vector(8 DOWNTO 0);
     L1619              :in std_logic_vector(8 DOWNTO 0);
     L1620              :in std_logic_vector(8 DOWNTO 0);
     L1621              :in std_logic_vector(8 DOWNTO 0);
     L1622              :in std_logic_vector(8 DOWNTO 0);
     L1623              :in std_logic_vector(8 DOWNTO 0);
     L1624              :in std_logic_vector(8 DOWNTO 0);
     L1625              :in std_logic_vector(8 DOWNTO 0);
     L1626              :in std_logic_vector(8 DOWNTO 0);
     L1627              :in std_logic_vector(8 DOWNTO 0);
     L1628              :in std_logic_vector(8 DOWNTO 0);
     L1629              :in std_logic_vector(8 DOWNTO 0);
     L1630              :in std_logic_vector(8 DOWNTO 0);
     L1631              :in std_logic_vector(8 DOWNTO 0);
     L1632              :in std_logic_vector(8 DOWNTO 0);
     L1633              :in std_logic_vector(8 DOWNTO 0);
     L1634              :in std_logic_vector(8 DOWNTO 0);
     L1635              :in std_logic_vector(8 DOWNTO 0);
     L1636              :in std_logic_vector(8 DOWNTO 0);
     L1637              :in std_logic_vector(8 DOWNTO 0);
     L1638              :in std_logic_vector(8 DOWNTO 0);
     L1639              :in std_logic_vector(8 DOWNTO 0);
     L1640              :in std_logic_vector(8 DOWNTO 0);
     L1641              :in std_logic_vector(8 DOWNTO 0);
     L1642              :in std_logic_vector(8 DOWNTO 0);
     L1643              :in std_logic_vector(8 DOWNTO 0);
     L1644              :in std_logic_vector(8 DOWNTO 0);
     L1645              :in std_logic_vector(8 DOWNTO 0);
     L1646              :in std_logic_vector(8 DOWNTO 0);
     L1647              :in std_logic_vector(8 DOWNTO 0);
     L1648              :in std_logic_vector(8 DOWNTO 0);
     L1649              :in std_logic_vector(8 DOWNTO 0);
     L1650              :in std_logic_vector(8 DOWNTO 0);
     L1651              :in std_logic_vector(8 DOWNTO 0);
     L1652              :in std_logic_vector(8 DOWNTO 0);
     L1653              :in std_logic_vector(8 DOWNTO 0);
     L1654              :in std_logic_vector(8 DOWNTO 0);
     L1655              :in std_logic_vector(8 DOWNTO 0);
     L1656              :in std_logic_vector(8 DOWNTO 0);
     L1657              :in std_logic_vector(8 DOWNTO 0);
     L1658              :in std_logic_vector(8 DOWNTO 0);
     L1659              :in std_logic_vector(8 DOWNTO 0);
     L1660              :in std_logic_vector(8 DOWNTO 0);
     L1661              :in std_logic_vector(8 DOWNTO 0);
     L1662              :in std_logic_vector(8 DOWNTO 0);
     L1663              :in std_logic_vector(8 DOWNTO 0);
     L1664              :in std_logic_vector(8 DOWNTO 0);
     L1665              :in std_logic_vector(8 DOWNTO 0);
     L1666              :in std_logic_vector(8 DOWNTO 0);
     L1667              :in std_logic_vector(8 DOWNTO 0);
     L1668              :in std_logic_vector(8 DOWNTO 0);
     L1669              :in std_logic_vector(8 DOWNTO 0);
     L1670              :in std_logic_vector(8 DOWNTO 0);
     L1671              :in std_logic_vector(8 DOWNTO 0);
     L1672              :in std_logic_vector(8 DOWNTO 0);
     L1673              :in std_logic_vector(8 DOWNTO 0);
     L1674              :in std_logic_vector(8 DOWNTO 0);
     L1675              :in std_logic_vector(8 DOWNTO 0);
     L1676              :in std_logic_vector(8 DOWNTO 0);
     L1677              :in std_logic_vector(8 DOWNTO 0);
     L1678              :in std_logic_vector(8 DOWNTO 0);
     L1679              :in std_logic_vector(8 DOWNTO 0);
     L1680              :in std_logic_vector(8 DOWNTO 0);
     L1681              :in std_logic_vector(8 DOWNTO 0);
     L1682              :in std_logic_vector(8 DOWNTO 0);
     L1683              :in std_logic_vector(8 DOWNTO 0);
     L1684              :in std_logic_vector(8 DOWNTO 0);
     L1685              :in std_logic_vector(8 DOWNTO 0);
     L1686              :in std_logic_vector(8 DOWNTO 0);
     L1687              :in std_logic_vector(8 DOWNTO 0);
     L1688              :in std_logic_vector(8 DOWNTO 0);
     L1689              :in std_logic_vector(8 DOWNTO 0);
     L1690              :in std_logic_vector(8 DOWNTO 0);
     L1691              :in std_logic_vector(8 DOWNTO 0);
     L1692              :in std_logic_vector(8 DOWNTO 0);
     L1693              :in std_logic_vector(8 DOWNTO 0);
     L1694              :in std_logic_vector(8 DOWNTO 0);
     L1695              :in std_logic_vector(8 DOWNTO 0);
     L1696              :in std_logic_vector(8 DOWNTO 0);
     L1697              :in std_logic_vector(8 DOWNTO 0);
     L1698              :in std_logic_vector(8 DOWNTO 0);
     L1699              :in std_logic_vector(8 DOWNTO 0);
     L1700              :in std_logic_vector(8 DOWNTO 0);
     L1701              :in std_logic_vector(8 DOWNTO 0);
     L1702              :in std_logic_vector(8 DOWNTO 0);
     L1703              :in std_logic_vector(8 DOWNTO 0);
     L1704              :in std_logic_vector(8 DOWNTO 0);
     L1705              :in std_logic_vector(8 DOWNTO 0);
     L1706              :in std_logic_vector(8 DOWNTO 0);
     L1707              :in std_logic_vector(8 DOWNTO 0);
     L1708              :in std_logic_vector(8 DOWNTO 0);
     L1709              :in std_logic_vector(8 DOWNTO 0);
     L1710              :in std_logic_vector(8 DOWNTO 0);
     L1711              :in std_logic_vector(8 DOWNTO 0);
     L1712              :in std_logic_vector(8 DOWNTO 0);
     L1713              :in std_logic_vector(8 DOWNTO 0);
     L1714              :in std_logic_vector(8 DOWNTO 0);
     L1715              :in std_logic_vector(8 DOWNTO 0);
     L1716              :in std_logic_vector(8 DOWNTO 0);
     L1717              :in std_logic_vector(8 DOWNTO 0);
     L1718              :in std_logic_vector(8 DOWNTO 0);
     L1719              :in std_logic_vector(8 DOWNTO 0);
     L1720              :in std_logic_vector(8 DOWNTO 0);
     L1721              :in std_logic_vector(8 DOWNTO 0);
     L1722              :in std_logic_vector(8 DOWNTO 0);
     L1723              :in std_logic_vector(8 DOWNTO 0);
     L1724              :in std_logic_vector(8 DOWNTO 0);
     L1725              :in std_logic_vector(8 DOWNTO 0);
     L1726              :in std_logic_vector(8 DOWNTO 0);
     L1727              :in std_logic_vector(8 DOWNTO 0);
     L1728              :in std_logic_vector(8 DOWNTO 0);
     L1729              :in std_logic_vector(8 DOWNTO 0);
     L1730              :in std_logic_vector(8 DOWNTO 0);
     L1731              :in std_logic_vector(8 DOWNTO 0);
     L1732              :in std_logic_vector(8 DOWNTO 0);
     L1733              :in std_logic_vector(8 DOWNTO 0);
     L1734              :in std_logic_vector(8 DOWNTO 0);
     L1735              :in std_logic_vector(8 DOWNTO 0);
     L1736              :in std_logic_vector(8 DOWNTO 0);
     L1737              :in std_logic_vector(8 DOWNTO 0);
     L1738              :in std_logic_vector(8 DOWNTO 0);
     L1739              :in std_logic_vector(8 DOWNTO 0);
     L1740              :in std_logic_vector(8 DOWNTO 0);
     L1741              :in std_logic_vector(8 DOWNTO 0);
     L1742              :in std_logic_vector(8 DOWNTO 0);
     L1743              :in std_logic_vector(8 DOWNTO 0);
     L1744              :in std_logic_vector(8 DOWNTO 0);
     L1745              :in std_logic_vector(8 DOWNTO 0);
     L1746              :in std_logic_vector(8 DOWNTO 0);
     L1747              :in std_logic_vector(8 DOWNTO 0);
     L1748              :in std_logic_vector(8 DOWNTO 0);
     L1749              :in std_logic_vector(8 DOWNTO 0);
     L1750              :in std_logic_vector(8 DOWNTO 0);
     L1751              :in std_logic_vector(8 DOWNTO 0);
     L1752              :in std_logic_vector(8 DOWNTO 0);
     L1753              :in std_logic_vector(8 DOWNTO 0);
     L1754              :in std_logic_vector(8 DOWNTO 0);
     L1755              :in std_logic_vector(8 DOWNTO 0);
     L1756              :in std_logic_vector(8 DOWNTO 0);
     L1757              :in std_logic_vector(8 DOWNTO 0);
     L1758              :in std_logic_vector(8 DOWNTO 0);
     L1759              :in std_logic_vector(8 DOWNTO 0);
     L1760              :in std_logic_vector(8 DOWNTO 0);
     L1761              :in std_logic_vector(8 DOWNTO 0);
     L1762              :in std_logic_vector(8 DOWNTO 0);
     L1763              :in std_logic_vector(8 DOWNTO 0);
     L1764              :in std_logic_vector(8 DOWNTO 0);
     L1765              :in std_logic_vector(8 DOWNTO 0);
     L1766              :in std_logic_vector(8 DOWNTO 0);
     L1767              :in std_logic_vector(8 DOWNTO 0);
     L1768              :in std_logic_vector(8 DOWNTO 0);
     L1769              :in std_logic_vector(8 DOWNTO 0);
     L1770              :in std_logic_vector(8 DOWNTO 0);
     L1771              :in std_logic_vector(8 DOWNTO 0);
     L1772              :in std_logic_vector(8 DOWNTO 0);
     L1773              :in std_logic_vector(8 DOWNTO 0);
     L1774              :in std_logic_vector(8 DOWNTO 0);
     L1775              :in std_logic_vector(8 DOWNTO 0);
     L1776              :in std_logic_vector(8 DOWNTO 0);
     L1777              :in std_logic_vector(8 DOWNTO 0);
     L1778              :in std_logic_vector(8 DOWNTO 0);
     L1779              :in std_logic_vector(8 DOWNTO 0);
     L1780              :in std_logic_vector(8 DOWNTO 0);
     L1781              :in std_logic_vector(8 DOWNTO 0);
     L1782              :in std_logic_vector(8 DOWNTO 0);
     L1783              :in std_logic_vector(8 DOWNTO 0);
     L1784              :in std_logic_vector(8 DOWNTO 0);
     L1785              :in std_logic_vector(8 DOWNTO 0);
     L1786              :in std_logic_vector(8 DOWNTO 0);
     L1787              :in std_logic_vector(8 DOWNTO 0);
     L1788              :in std_logic_vector(8 DOWNTO 0);
     L1789              :in std_logic_vector(8 DOWNTO 0);
     L1790              :in std_logic_vector(8 DOWNTO 0);
     L1791              :in std_logic_vector(8 DOWNTO 0);
     L1792              :in std_logic_vector(8 DOWNTO 0);
     L1793              :in std_logic_vector(8 DOWNTO 0);
     L1794              :in std_logic_vector(8 DOWNTO 0);
     L1795              :in std_logic_vector(8 DOWNTO 0);
     L1796              :in std_logic_vector(8 DOWNTO 0);
     L1797              :in std_logic_vector(8 DOWNTO 0);
     L1798              :in std_logic_vector(8 DOWNTO 0);
     L1799              :in std_logic_vector(8 DOWNTO 0);
     L1800              :in std_logic_vector(8 DOWNTO 0);
     L1801              :in std_logic_vector(8 DOWNTO 0);
     L1802              :in std_logic_vector(8 DOWNTO 0);
     L1803              :in std_logic_vector(8 DOWNTO 0);
     L1804              :in std_logic_vector(8 DOWNTO 0);
     L1805              :in std_logic_vector(8 DOWNTO 0);
     L1806              :in std_logic_vector(8 DOWNTO 0);
     L1807              :in std_logic_vector(8 DOWNTO 0);
     L1808              :in std_logic_vector(8 DOWNTO 0);
     L1809              :in std_logic_vector(8 DOWNTO 0);
     L1810              :in std_logic_vector(8 DOWNTO 0);
     L1811              :in std_logic_vector(8 DOWNTO 0);
     L1812              :in std_logic_vector(8 DOWNTO 0);
     L1813              :in std_logic_vector(8 DOWNTO 0);
     L1814              :in std_logic_vector(8 DOWNTO 0);
     L1815              :in std_logic_vector(8 DOWNTO 0);
     L1816              :in std_logic_vector(8 DOWNTO 0);
     L1817              :in std_logic_vector(8 DOWNTO 0);
     L1818              :in std_logic_vector(8 DOWNTO 0);
     L1819              :in std_logic_vector(8 DOWNTO 0);
     L1820              :in std_logic_vector(8 DOWNTO 0);
     L1821              :in std_logic_vector(8 DOWNTO 0);
     L1822              :in std_logic_vector(8 DOWNTO 0);
     L1823              :in std_logic_vector(8 DOWNTO 0);
     L1824              :in std_logic_vector(8 DOWNTO 0);
     L1825              :in std_logic_vector(8 DOWNTO 0);
     L1826              :in std_logic_vector(8 DOWNTO 0);
     L1827              :in std_logic_vector(8 DOWNTO 0);
     L1828              :in std_logic_vector(8 DOWNTO 0);
     L1829              :in std_logic_vector(8 DOWNTO 0);
     L1830              :in std_logic_vector(8 DOWNTO 0);
     L1831              :in std_logic_vector(8 DOWNTO 0);
     L1832              :in std_logic_vector(8 DOWNTO 0);
     L1833              :in std_logic_vector(8 DOWNTO 0);
     L1834              :in std_logic_vector(8 DOWNTO 0);
     L1835              :in std_logic_vector(8 DOWNTO 0);
     L1836              :in std_logic_vector(8 DOWNTO 0);
     L1837              :in std_logic_vector(8 DOWNTO 0);
     L1838              :in std_logic_vector(8 DOWNTO 0);
     L1839              :in std_logic_vector(8 DOWNTO 0);
     L1840              :in std_logic_vector(8 DOWNTO 0);
     L1841              :in std_logic_vector(8 DOWNTO 0);
     L1842              :in std_logic_vector(8 DOWNTO 0);
     L1843              :in std_logic_vector(8 DOWNTO 0);
     L1844              :in std_logic_vector(8 DOWNTO 0);
     L1845              :in std_logic_vector(8 DOWNTO 0);
     L1846              :in std_logic_vector(8 DOWNTO 0);
     L1847              :in std_logic_vector(8 DOWNTO 0);
     L1848              :in std_logic_vector(8 DOWNTO 0);
     L1849              :in std_logic_vector(8 DOWNTO 0);
     L1850              :in std_logic_vector(8 DOWNTO 0);
     L1851              :in std_logic_vector(8 DOWNTO 0);
     L1852              :in std_logic_vector(8 DOWNTO 0);
     L1853              :in std_logic_vector(8 DOWNTO 0);
     L1854              :in std_logic_vector(8 DOWNTO 0);
     L1855              :in std_logic_vector(8 DOWNTO 0);
     L1856              :in std_logic_vector(8 DOWNTO 0);
     L1857              :in std_logic_vector(8 DOWNTO 0);
     L1858              :in std_logic_vector(8 DOWNTO 0);
     L1859              :in std_logic_vector(8 DOWNTO 0);
     L1860              :in std_logic_vector(8 DOWNTO 0);
     L1861              :in std_logic_vector(8 DOWNTO 0);
     L1862              :in std_logic_vector(8 DOWNTO 0);
     L1863              :in std_logic_vector(8 DOWNTO 0);
     L1864              :in std_logic_vector(8 DOWNTO 0);
     L1865              :in std_logic_vector(8 DOWNTO 0);
     L1866              :in std_logic_vector(8 DOWNTO 0);
     L1867              :in std_logic_vector(8 DOWNTO 0);
     L1868              :in std_logic_vector(8 DOWNTO 0);
     L1869              :in std_logic_vector(8 DOWNTO 0);
     L1870              :in std_logic_vector(8 DOWNTO 0);
     L1871              :in std_logic_vector(8 DOWNTO 0);
     L1872              :in std_logic_vector(8 DOWNTO 0);
     L1873              :in std_logic_vector(8 DOWNTO 0);
     L1874              :in std_logic_vector(8 DOWNTO 0);
     L1875              :in std_logic_vector(8 DOWNTO 0);
     L1876              :in std_logic_vector(8 DOWNTO 0);
     L1877              :in std_logic_vector(8 DOWNTO 0);
     L1878              :in std_logic_vector(8 DOWNTO 0);
     L1879              :in std_logic_vector(8 DOWNTO 0);
     L1880              :in std_logic_vector(8 DOWNTO 0);
     L1881              :in std_logic_vector(8 DOWNTO 0);
     L1882              :in std_logic_vector(8 DOWNTO 0);
     L1883              :in std_logic_vector(8 DOWNTO 0);
     L1884              :in std_logic_vector(8 DOWNTO 0);
     L1885              :in std_logic_vector(8 DOWNTO 0);
     L1886              :in std_logic_vector(8 DOWNTO 0);
     L1887              :in std_logic_vector(8 DOWNTO 0);
     L1888              :in std_logic_vector(8 DOWNTO 0);
     L1889              :in std_logic_vector(8 DOWNTO 0);
     L1890              :in std_logic_vector(8 DOWNTO 0);
     L1891              :in std_logic_vector(8 DOWNTO 0);
     L1892              :in std_logic_vector(8 DOWNTO 0);
     L1893              :in std_logic_vector(8 DOWNTO 0);
     L1894              :in std_logic_vector(8 DOWNTO 0);
     L1895              :in std_logic_vector(8 DOWNTO 0);
     L1896              :in std_logic_vector(8 DOWNTO 0);
     L1897              :in std_logic_vector(8 DOWNTO 0);
     L1898              :in std_logic_vector(8 DOWNTO 0);
     L1899              :in std_logic_vector(8 DOWNTO 0);
     L1900              :in std_logic_vector(8 DOWNTO 0);
     L1901              :in std_logic_vector(8 DOWNTO 0);
     L1902              :in std_logic_vector(8 DOWNTO 0);
     L1903              :in std_logic_vector(8 DOWNTO 0);
     L1904              :in std_logic_vector(8 DOWNTO 0);
     L1905              :in std_logic_vector(8 DOWNTO 0);
     L1906              :in std_logic_vector(8 DOWNTO 0);
     L1907              :in std_logic_vector(8 DOWNTO 0);
     L1908              :in std_logic_vector(8 DOWNTO 0);
     L1909              :in std_logic_vector(8 DOWNTO 0);
     L1910              :in std_logic_vector(8 DOWNTO 0);
     L1911              :in std_logic_vector(8 DOWNTO 0);
     L1912              :in std_logic_vector(8 DOWNTO 0);
     L1913              :in std_logic_vector(8 DOWNTO 0);
     L1914              :in std_logic_vector(8 DOWNTO 0);
     L1915              :in std_logic_vector(8 DOWNTO 0);
     L1916              :in std_logic_vector(8 DOWNTO 0);
     L1917              :in std_logic_vector(8 DOWNTO 0);
     L1918              :in std_logic_vector(8 DOWNTO 0);
     L1919              :in std_logic_vector(8 DOWNTO 0);
     L1920              :in std_logic_vector(8 DOWNTO 0);
     L1921              :in std_logic_vector(8 DOWNTO 0);
     L1922              :in std_logic_vector(8 DOWNTO 0);
     L1923              :in std_logic_vector(8 DOWNTO 0);
     L1924              :in std_logic_vector(8 DOWNTO 0);
     L1925              :in std_logic_vector(8 DOWNTO 0);
     L1926              :in std_logic_vector(8 DOWNTO 0);
     L1927              :in std_logic_vector(8 DOWNTO 0);
     L1928              :in std_logic_vector(8 DOWNTO 0);
     L1929              :in std_logic_vector(8 DOWNTO 0);
     L1930              :in std_logic_vector(8 DOWNTO 0);
     L1931              :in std_logic_vector(8 DOWNTO 0);
     L1932              :in std_logic_vector(8 DOWNTO 0);
     L1933              :in std_logic_vector(8 DOWNTO 0);
     L1934              :in std_logic_vector(8 DOWNTO 0);
     L1935              :in std_logic_vector(8 DOWNTO 0);
     L1936              :in std_logic_vector(8 DOWNTO 0);
     L1937              :in std_logic_vector(8 DOWNTO 0);
     L1938              :in std_logic_vector(8 DOWNTO 0);
     L1939              :in std_logic_vector(8 DOWNTO 0);
     L1940              :in std_logic_vector(8 DOWNTO 0);
     L1941              :in std_logic_vector(8 DOWNTO 0);
     L1942              :in std_logic_vector(8 DOWNTO 0);
     L1943              :in std_logic_vector(8 DOWNTO 0);
     L1944              :in std_logic_vector(8 DOWNTO 0);
     L1945              :in std_logic_vector(8 DOWNTO 0);
     L1946              :in std_logic_vector(8 DOWNTO 0);
     L1947              :in std_logic_vector(8 DOWNTO 0);
     L1948              :in std_logic_vector(8 DOWNTO 0);
     L1949              :in std_logic_vector(8 DOWNTO 0);
     L1950              :in std_logic_vector(8 DOWNTO 0);
     L1951              :in std_logic_vector(8 DOWNTO 0);
     L1952              :in std_logic_vector(8 DOWNTO 0);
     L1953              :in std_logic_vector(8 DOWNTO 0);
     L1954              :in std_logic_vector(8 DOWNTO 0);
     L1955              :in std_logic_vector(8 DOWNTO 0);
     L1956              :in std_logic_vector(8 DOWNTO 0);
     L1957              :in std_logic_vector(8 DOWNTO 0);
     L1958              :in std_logic_vector(8 DOWNTO 0);
     L1959              :in std_logic_vector(8 DOWNTO 0);
     L1960              :in std_logic_vector(8 DOWNTO 0);
     L1961              :in std_logic_vector(8 DOWNTO 0);
     L1962              :in std_logic_vector(8 DOWNTO 0);
     L1963              :in std_logic_vector(8 DOWNTO 0);
     L1964              :in std_logic_vector(8 DOWNTO 0);
     L1965              :in std_logic_vector(8 DOWNTO 0);
     L1966              :in std_logic_vector(8 DOWNTO 0);
     L1967              :in std_logic_vector(8 DOWNTO 0);
     L1968              :in std_logic_vector(8 DOWNTO 0);
     L1969              :in std_logic_vector(8 DOWNTO 0);
     L1970              :in std_logic_vector(8 DOWNTO 0);
     L1971              :in std_logic_vector(8 DOWNTO 0);
     L1972              :in std_logic_vector(8 DOWNTO 0);
     L1973              :in std_logic_vector(8 DOWNTO 0);
     L1974              :in std_logic_vector(8 DOWNTO 0);
     L1975              :in std_logic_vector(8 DOWNTO 0);
     L1976              :in std_logic_vector(8 DOWNTO 0);
     L1977              :in std_logic_vector(8 DOWNTO 0);
     L1978              :in std_logic_vector(8 DOWNTO 0);
     L1979              :in std_logic_vector(8 DOWNTO 0);
     L1980              :in std_logic_vector(8 DOWNTO 0);
     L1981              :in std_logic_vector(8 DOWNTO 0);
     L1982              :in std_logic_vector(8 DOWNTO 0);
     L1983              :in std_logic_vector(8 DOWNTO 0);
     L1984              :in std_logic_vector(8 DOWNTO 0);
     L1985              :in std_logic_vector(8 DOWNTO 0);
     L1986              :in std_logic_vector(8 DOWNTO 0);
     L1987              :in std_logic_vector(8 DOWNTO 0);
     L1988              :in std_logic_vector(8 DOWNTO 0);
     L1989              :in std_logic_vector(8 DOWNTO 0);
     L1990              :in std_logic_vector(8 DOWNTO 0);
     L1991              :in std_logic_vector(8 DOWNTO 0);
     L1992              :in std_logic_vector(8 DOWNTO 0);
     L1993              :in std_logic_vector(8 DOWNTO 0);
     L1994              :in std_logic_vector(8 DOWNTO 0);
     L1995              :in std_logic_vector(8 DOWNTO 0);
     L1996              :in std_logic_vector(8 DOWNTO 0);
     L1997              :in std_logic_vector(8 DOWNTO 0);
     L1998              :in std_logic_vector(8 DOWNTO 0);
     L1999              :in std_logic_vector(8 DOWNTO 0);
     L2000              :in std_logic_vector(8 DOWNTO 0);
     L2001              :in std_logic_vector(8 DOWNTO 0);
     L2002              :in std_logic_vector(8 DOWNTO 0);
     L2003              :in std_logic_vector(8 DOWNTO 0);
     L2004              :in std_logic_vector(8 DOWNTO 0);
     L2005              :in std_logic_vector(8 DOWNTO 0);
     L2006              :in std_logic_vector(8 DOWNTO 0);
     L2007              :in std_logic_vector(8 DOWNTO 0);
     L2008              :in std_logic_vector(8 DOWNTO 0);
     L2009              :in std_logic_vector(8 DOWNTO 0);
     L2010              :in std_logic_vector(8 DOWNTO 0);
     L2011              :in std_logic_vector(8 DOWNTO 0);
     L2012              :in std_logic_vector(8 DOWNTO 0);
     L2013              :in std_logic_vector(8 DOWNTO 0);
     L2014              :in std_logic_vector(8 DOWNTO 0);
     L2015              :in std_logic_vector(8 DOWNTO 0);
     L2016              :in std_logic_vector(8 DOWNTO 0);
     L2017              :in std_logic_vector(8 DOWNTO 0);
     L2018              :in std_logic_vector(8 DOWNTO 0);
     L2019              :in std_logic_vector(8 DOWNTO 0);
     L2020              :in std_logic_vector(8 DOWNTO 0);
     L2021              :in std_logic_vector(8 DOWNTO 0);
     L2022              :in std_logic_vector(8 DOWNTO 0);
     L2023              :in std_logic_vector(8 DOWNTO 0);
     L2024              :in std_logic_vector(8 DOWNTO 0);
     L2025              :in std_logic_vector(8 DOWNTO 0);
     L2026              :in std_logic_vector(8 DOWNTO 0);
     L2027              :in std_logic_vector(8 DOWNTO 0);
     L2028              :in std_logic_vector(8 DOWNTO 0);
     L2029              :in std_logic_vector(8 DOWNTO 0);
     L2030              :in std_logic_vector(8 DOWNTO 0);
     L2031              :in std_logic_vector(8 DOWNTO 0);
     L2032              :in std_logic_vector(8 DOWNTO 0);
     L2033              :in std_logic_vector(8 DOWNTO 0);
     L2034              :in std_logic_vector(8 DOWNTO 0);
     L2035              :in std_logic_vector(8 DOWNTO 0);
     L2036              :in std_logic_vector(8 DOWNTO 0);
     L2037              :in std_logic_vector(8 DOWNTO 0);
     L2038              :in std_logic_vector(8 DOWNTO 0);
     L2039              :in std_logic_vector(8 DOWNTO 0);
     L2040              :in std_logic_vector(8 DOWNTO 0);
     L2041              :in std_logic_vector(8 DOWNTO 0);
     L2042              :in std_logic_vector(8 DOWNTO 0);
     L2043              :in std_logic_vector(8 DOWNTO 0);
     L2044              :in std_logic_vector(8 DOWNTO 0);
     L2045              :in std_logic_vector(8 DOWNTO 0);
     L2046              :in std_logic_vector(8 DOWNTO 0);
     L2047              :in std_logic_vector(8 DOWNTO 0);
     L2048              :in std_logic_vector(8 DOWNTO 0);
     L2049              :in std_logic_vector(8 DOWNTO 0);
     L2050              :in std_logic_vector(8 DOWNTO 0);
     L2051              :in std_logic_vector(8 DOWNTO 0);
     L2052              :in std_logic_vector(8 DOWNTO 0);
     L2053              :in std_logic_vector(8 DOWNTO 0);
     L2054              :in std_logic_vector(8 DOWNTO 0);
     L2055              :in std_logic_vector(8 DOWNTO 0);
     L2056              :in std_logic_vector(8 DOWNTO 0);
     L2057              :in std_logic_vector(8 DOWNTO 0);
     L2058              :in std_logic_vector(8 DOWNTO 0);
     L2059              :in std_logic_vector(8 DOWNTO 0);
     L2060              :in std_logic_vector(8 DOWNTO 0);
     L2061              :in std_logic_vector(8 DOWNTO 0);
     L2062              :in std_logic_vector(8 DOWNTO 0);
     L2063              :in std_logic_vector(8 DOWNTO 0);
     L2064              :in std_logic_vector(8 DOWNTO 0);
     L2065              :in std_logic_vector(8 DOWNTO 0);
     L2066              :in std_logic_vector(8 DOWNTO 0);
     L2067              :in std_logic_vector(8 DOWNTO 0);
     L2068              :in std_logic_vector(8 DOWNTO 0);
     L2069              :in std_logic_vector(8 DOWNTO 0);
     L2070              :in std_logic_vector(8 DOWNTO 0);
     L2071              :in std_logic_vector(8 DOWNTO 0);
     L2072              :in std_logic_vector(8 DOWNTO 0);
     L2073              :in std_logic_vector(8 DOWNTO 0);
     L2074              :in std_logic_vector(8 DOWNTO 0);
     L2075              :in std_logic_vector(8 DOWNTO 0);
     L2076              :in std_logic_vector(8 DOWNTO 0);
     L2077              :in std_logic_vector(8 DOWNTO 0);
     L2078              :in std_logic_vector(8 DOWNTO 0);
     L2079              :in std_logic_vector(8 DOWNTO 0);
     L2080              :in std_logic_vector(8 DOWNTO 0);
     L2081              :in std_logic_vector(8 DOWNTO 0);
     L2082              :in std_logic_vector(8 DOWNTO 0);
     L2083              :in std_logic_vector(8 DOWNTO 0);
     L2084              :in std_logic_vector(8 DOWNTO 0);
     L2085              :in std_logic_vector(8 DOWNTO 0);
     L2086              :in std_logic_vector(8 DOWNTO 0);
     L2087              :in std_logic_vector(8 DOWNTO 0);
     L2088              :in std_logic_vector(8 DOWNTO 0);
     L2089              :in std_logic_vector(8 DOWNTO 0);
     L2090              :in std_logic_vector(8 DOWNTO 0);
     L2091              :in std_logic_vector(8 DOWNTO 0);
     L2092              :in std_logic_vector(8 DOWNTO 0);
     L2093              :in std_logic_vector(8 DOWNTO 0);
     L2094              :in std_logic_vector(8 DOWNTO 0);
     L2095              :in std_logic_vector(8 DOWNTO 0);
     L2096              :in std_logic_vector(8 DOWNTO 0);
     L2097              :in std_logic_vector(8 DOWNTO 0);
     L2098              :in std_logic_vector(8 DOWNTO 0);
     L2099              :in std_logic_vector(8 DOWNTO 0);
     L2100              :in std_logic_vector(8 DOWNTO 0);
     L2101              :in std_logic_vector(8 DOWNTO 0);
     L2102              :in std_logic_vector(8 DOWNTO 0);
     L2103              :in std_logic_vector(8 DOWNTO 0);
     L2104              :in std_logic_vector(8 DOWNTO 0);
     L2105              :in std_logic_vector(8 DOWNTO 0);
     L2106              :in std_logic_vector(8 DOWNTO 0);
     L2107              :in std_logic_vector(8 DOWNTO 0);
     L2108              :in std_logic_vector(8 DOWNTO 0);
     L2109              :in std_logic_vector(8 DOWNTO 0);
     L2110              :in std_logic_vector(8 DOWNTO 0);
     L2111              :in std_logic_vector(8 DOWNTO 0);
     L2112              :in std_logic_vector(8 DOWNTO 0);
     L2113              :in std_logic_vector(8 DOWNTO 0);
     L2114              :in std_logic_vector(8 DOWNTO 0);
     L2115              :in std_logic_vector(8 DOWNTO 0);
     L2116              :in std_logic_vector(8 DOWNTO 0);
     L2117              :in std_logic_vector(8 DOWNTO 0);
     L2118              :in std_logic_vector(8 DOWNTO 0);
     L2119              :in std_logic_vector(8 DOWNTO 0);
     L2120              :in std_logic_vector(8 DOWNTO 0);
     L2121              :in std_logic_vector(8 DOWNTO 0);
     L2122              :in std_logic_vector(8 DOWNTO 0);
     L2123              :in std_logic_vector(8 DOWNTO 0);
     L2124              :in std_logic_vector(8 DOWNTO 0);
     L2125              :in std_logic_vector(8 DOWNTO 0);
     L2126              :in std_logic_vector(8 DOWNTO 0);
     L2127              :in std_logic_vector(8 DOWNTO 0);
     L2128              :in std_logic_vector(8 DOWNTO 0);
     L2129              :in std_logic_vector(8 DOWNTO 0);
     L2130              :in std_logic_vector(8 DOWNTO 0);
     L2131              :in std_logic_vector(8 DOWNTO 0);
     L2132              :in std_logic_vector(8 DOWNTO 0);
     L2133              :in std_logic_vector(8 DOWNTO 0);
     L2134              :in std_logic_vector(8 DOWNTO 0);
     L2135              :in std_logic_vector(8 DOWNTO 0);
     L2136              :in std_logic_vector(8 DOWNTO 0);
     L2137              :in std_logic_vector(8 DOWNTO 0);
     L2138              :in std_logic_vector(8 DOWNTO 0);
     L2139              :in std_logic_vector(8 DOWNTO 0);
     L2140              :in std_logic_vector(8 DOWNTO 0);
     L2141              :in std_logic_vector(8 DOWNTO 0);
     L2142              :in std_logic_vector(8 DOWNTO 0);
     L2143              :in std_logic_vector(8 DOWNTO 0);
     L2144              :in std_logic_vector(8 DOWNTO 0);
     L2145              :in std_logic_vector(8 DOWNTO 0);
     L2146              :in std_logic_vector(8 DOWNTO 0);
     L2147              :in std_logic_vector(8 DOWNTO 0);
     L2148              :in std_logic_vector(8 DOWNTO 0);
     L2149              :in std_logic_vector(8 DOWNTO 0);
     L2150              :in std_logic_vector(8 DOWNTO 0);
     L2151              :in std_logic_vector(8 DOWNTO 0);
     L2152              :in std_logic_vector(8 DOWNTO 0);
     L2153              :in std_logic_vector(8 DOWNTO 0);
     L2154              :in std_logic_vector(8 DOWNTO 0);
     L2155              :in std_logic_vector(8 DOWNTO 0);
     L2156              :in std_logic_vector(8 DOWNTO 0);
     L2157              :in std_logic_vector(8 DOWNTO 0);
     L2158              :in std_logic_vector(8 DOWNTO 0);
     L2159              :in std_logic_vector(8 DOWNTO 0);
     L2160              :in std_logic_vector(8 DOWNTO 0);
     L2161              :in std_logic_vector(8 DOWNTO 0);
     L2162              :in std_logic_vector(8 DOWNTO 0);
     L2163              :in std_logic_vector(8 DOWNTO 0);
     L2164              :in std_logic_vector(8 DOWNTO 0);
     L2165              :in std_logic_vector(8 DOWNTO 0);
     L2166              :in std_logic_vector(8 DOWNTO 0);
     L2167              :in std_logic_vector(8 DOWNTO 0);
     L2168              :in std_logic_vector(8 DOWNTO 0);
     L2169              :in std_logic_vector(8 DOWNTO 0);
     L2170              :in std_logic_vector(8 DOWNTO 0);
     L2171              :in std_logic_vector(8 DOWNTO 0);
     L2172              :in std_logic_vector(8 DOWNTO 0);
     L2173              :in std_logic_vector(8 DOWNTO 0);
     L2174              :in std_logic_vector(8 DOWNTO 0);
     L2175              :in std_logic_vector(8 DOWNTO 0);
     L2176              :in std_logic_vector(8 DOWNTO 0);
     L2177              :in std_logic_vector(8 DOWNTO 0);
     L2178              :in std_logic_vector(8 DOWNTO 0);
     L2179              :in std_logic_vector(8 DOWNTO 0);
     L2180              :in std_logic_vector(8 DOWNTO 0);
     L2181              :in std_logic_vector(8 DOWNTO 0);
     L2182              :in std_logic_vector(8 DOWNTO 0);
     L2183              :in std_logic_vector(8 DOWNTO 0);
     L2184              :in std_logic_vector(8 DOWNTO 0);
     L2185              :in std_logic_vector(8 DOWNTO 0);
     L2186              :in std_logic_vector(8 DOWNTO 0);
     L2187              :in std_logic_vector(8 DOWNTO 0);
     L2188              :in std_logic_vector(8 DOWNTO 0);
     L2189              :in std_logic_vector(8 DOWNTO 0);
     L2190              :in std_logic_vector(8 DOWNTO 0);
     L2191              :in std_logic_vector(8 DOWNTO 0);
     L2192              :in std_logic_vector(8 DOWNTO 0);
     L2193              :in std_logic_vector(8 DOWNTO 0);
     L2194              :in std_logic_vector(8 DOWNTO 0);
     L2195              :in std_logic_vector(8 DOWNTO 0);
     L2196              :in std_logic_vector(8 DOWNTO 0);
     L2197              :in std_logic_vector(8 DOWNTO 0);
     L2198              :in std_logic_vector(8 DOWNTO 0);
     L2199              :in std_logic_vector(8 DOWNTO 0);
     L2200              :in std_logic_vector(8 DOWNTO 0);
     L2201              :in std_logic_vector(8 DOWNTO 0);
     L2202              :in std_logic_vector(8 DOWNTO 0);
     L2203              :in std_logic_vector(8 DOWNTO 0);
     L2204              :in std_logic_vector(8 DOWNTO 0);
     L2205              :in std_logic_vector(8 DOWNTO 0);
     L2206              :in std_logic_vector(8 DOWNTO 0);
     L2207              :in std_logic_vector(8 DOWNTO 0);
     L2208              :in std_logic_vector(8 DOWNTO 0);
     L2209              :in std_logic_vector(8 DOWNTO 0);
     L2210              :in std_logic_vector(8 DOWNTO 0);
     L2211              :in std_logic_vector(8 DOWNTO 0);
     L2212              :in std_logic_vector(8 DOWNTO 0);
     L2213              :in std_logic_vector(8 DOWNTO 0);
     L2214              :in std_logic_vector(8 DOWNTO 0);
     L2215              :in std_logic_vector(8 DOWNTO 0);
     L2216              :in std_logic_vector(8 DOWNTO 0);
     L2217              :in std_logic_vector(8 DOWNTO 0);
     L2218              :in std_logic_vector(8 DOWNTO 0);
     L2219              :in std_logic_vector(8 DOWNTO 0);
     L2220              :in std_logic_vector(8 DOWNTO 0);
     L2221              :in std_logic_vector(8 DOWNTO 0);
     L2222              :in std_logic_vector(8 DOWNTO 0);
     L2223              :in std_logic_vector(8 DOWNTO 0);
     L2224              :in std_logic_vector(8 DOWNTO 0);
     L2225              :in std_logic_vector(8 DOWNTO 0);
     L2226              :in std_logic_vector(8 DOWNTO 0);
     L2227              :in std_logic_vector(8 DOWNTO 0);
     L2228              :in std_logic_vector(8 DOWNTO 0);
     L2229              :in std_logic_vector(8 DOWNTO 0);
     L2230              :in std_logic_vector(8 DOWNTO 0);
     L2231              :in std_logic_vector(8 DOWNTO 0);
     L2232              :in std_logic_vector(8 DOWNTO 0);
     L2233              :in std_logic_vector(8 DOWNTO 0);
     L2234              :in std_logic_vector(8 DOWNTO 0);
     L2235              :in std_logic_vector(8 DOWNTO 0);
     L2236              :in std_logic_vector(8 DOWNTO 0);
     L2237              :in std_logic_vector(8 DOWNTO 0);
     L2238              :in std_logic_vector(8 DOWNTO 0);
     L2239              :in std_logic_vector(8 DOWNTO 0);
     L2240              :in std_logic_vector(8 DOWNTO 0);
     L2241              :in std_logic_vector(8 DOWNTO 0);
     L2242              :in std_logic_vector(8 DOWNTO 0);
     L2243              :in std_logic_vector(8 DOWNTO 0);
     L2244              :in std_logic_vector(8 DOWNTO 0);
     L2245              :in std_logic_vector(8 DOWNTO 0);
     L2246              :in std_logic_vector(8 DOWNTO 0);
     L2247              :in std_logic_vector(8 DOWNTO 0);
     L2248              :in std_logic_vector(8 DOWNTO 0);
     L2249              :in std_logic_vector(8 DOWNTO 0);
     L2250              :in std_logic_vector(8 DOWNTO 0);
     L2251              :in std_logic_vector(8 DOWNTO 0);
     L2252              :in std_logic_vector(8 DOWNTO 0);
     L2253              :in std_logic_vector(8 DOWNTO 0);
     L2254              :in std_logic_vector(8 DOWNTO 0);
     L2255              :in std_logic_vector(8 DOWNTO 0);
     L2256              :in std_logic_vector(8 DOWNTO 0);
     L2257              :in std_logic_vector(8 DOWNTO 0);
     L2258              :in std_logic_vector(8 DOWNTO 0);
     L2259              :in std_logic_vector(8 DOWNTO 0);
     L2260              :in std_logic_vector(8 DOWNTO 0);
     L2261              :in std_logic_vector(8 DOWNTO 0);
     L2262              :in std_logic_vector(8 DOWNTO 0);
     L2263              :in std_logic_vector(8 DOWNTO 0);
     L2264              :in std_logic_vector(8 DOWNTO 0);
     L2265              :in std_logic_vector(8 DOWNTO 0);
     L2266              :in std_logic_vector(8 DOWNTO 0);
     L2267              :in std_logic_vector(8 DOWNTO 0);
     L2268              :in std_logic_vector(8 DOWNTO 0);
     L2269              :in std_logic_vector(8 DOWNTO 0);
     L2270              :in std_logic_vector(8 DOWNTO 0);
     L2271              :in std_logic_vector(8 DOWNTO 0);
     L2272              :in std_logic_vector(8 DOWNTO 0);
     L2273              :in std_logic_vector(8 DOWNTO 0);
     L2274              :in std_logic_vector(8 DOWNTO 0);
     L2275              :in std_logic_vector(8 DOWNTO 0);
     L2276              :in std_logic_vector(8 DOWNTO 0);
     L2277              :in std_logic_vector(8 DOWNTO 0);
     L2278              :in std_logic_vector(8 DOWNTO 0);
     L2279              :in std_logic_vector(8 DOWNTO 0);
     L2280              :in std_logic_vector(8 DOWNTO 0);
     L2281              :in std_logic_vector(8 DOWNTO 0);
     L2282              :in std_logic_vector(8 DOWNTO 0);
     L2283              :in std_logic_vector(8 DOWNTO 0);
     L2284              :in std_logic_vector(8 DOWNTO 0);
     L2285              :in std_logic_vector(8 DOWNTO 0);
     L2286              :in std_logic_vector(8 DOWNTO 0);
     L2287              :in std_logic_vector(8 DOWNTO 0);
     L2288              :in std_logic_vector(8 DOWNTO 0);
     L2289              :in std_logic_vector(8 DOWNTO 0);
     L2290              :in std_logic_vector(8 DOWNTO 0);
     L2291              :in std_logic_vector(8 DOWNTO 0);
     L2292              :in std_logic_vector(8 DOWNTO 0);
     L2293              :in std_logic_vector(8 DOWNTO 0);
     L2294              :in std_logic_vector(8 DOWNTO 0);
     L2295              :in std_logic_vector(8 DOWNTO 0);
     L2296              :in std_logic_vector(8 DOWNTO 0);
     L2297              :in std_logic_vector(8 DOWNTO 0);
     L2298              :in std_logic_vector(8 DOWNTO 0);
     L2299              :in std_logic_vector(8 DOWNTO 0);
     L2300              :in std_logic_vector(8 DOWNTO 0);
     L2301              :in std_logic_vector(8 DOWNTO 0);
     L2302              :in std_logic_vector(8 DOWNTO 0);
     L2303              :in std_logic_vector(8 DOWNTO 0);
     L2304              :in std_logic_vector(8 DOWNTO 0);
     Z1            :out std_logic;
     Z2            :out std_logic;
     Z3            :out std_logic;
     Z4            :out std_logic;
     Z5            :out std_logic;
     Z6            :out std_logic;
     Z7            :out std_logic;
     Z8            :out std_logic;
     Z9            :out std_logic;
     Z10            :out std_logic;
     Z11            :out std_logic;
     Z12            :out std_logic;
     Z13            :out std_logic;
     Z14            :out std_logic;
     Z15            :out std_logic;
     Z16            :out std_logic;
     Z17            :out std_logic;
     Z18            :out std_logic;
     Z19            :out std_logic;
     Z20            :out std_logic;
     Z21            :out std_logic;
     Z22            :out std_logic;
     Z23            :out std_logic;
     Z24            :out std_logic;
     Z25            :out std_logic;
     Z26            :out std_logic;
     Z27            :out std_logic;
     Z28            :out std_logic;
     Z29            :out std_logic;
     Z30            :out std_logic;
     Z31            :out std_logic;
     Z32            :out std_logic;
     Z33            :out std_logic;
     Z34            :out std_logic;
     Z35            :out std_logic;
     Z36            :out std_logic;
     Z37            :out std_logic;
     Z38            :out std_logic;
     Z39            :out std_logic;
     Z40            :out std_logic;
     Z41            :out std_logic;
     Z42            :out std_logic;
     Z43            :out std_logic;
     Z44            :out std_logic;
     Z45            :out std_logic;
     Z46            :out std_logic;
     Z47            :out std_logic;
     Z48            :out std_logic;
     Z49            :out std_logic;
     Z50            :out std_logic;
     Z51            :out std_logic;
     Z52            :out std_logic;
     Z53            :out std_logic;
     Z54            :out std_logic;
     Z55            :out std_logic;
     Z56            :out std_logic;
     Z57            :out std_logic;
     Z58            :out std_logic;
     Z59            :out std_logic;
     Z60            :out std_logic;
     Z61            :out std_logic;
     Z62            :out std_logic;
     Z63            :out std_logic;
     Z64            :out std_logic;
     Z65            :out std_logic;
     Z66            :out std_logic;
     Z67            :out std_logic;
     Z68            :out std_logic;
     Z69            :out std_logic;
     Z70            :out std_logic;
     Z71            :out std_logic;
     Z72            :out std_logic;
     Z73            :out std_logic;
     Z74            :out std_logic;
     Z75            :out std_logic;
     Z76            :out std_logic;
     Z77            :out std_logic;
     Z78            :out std_logic;
     Z79            :out std_logic;
     Z80            :out std_logic;
     Z81            :out std_logic;
     Z82            :out std_logic;
     Z83            :out std_logic;
     Z84            :out std_logic;
     Z85            :out std_logic;
     Z86            :out std_logic;
     Z87            :out std_logic;
     Z88            :out std_logic;
     Z89            :out std_logic;
     Z90            :out std_logic;
     Z91            :out std_logic;
     Z92            :out std_logic;
     Z93            :out std_logic;
     Z94            :out std_logic;
     Z95            :out std_logic;
     Z96            :out std_logic;
     Z97            :out std_logic;
     Z98            :out std_logic;
     Z99            :out std_logic;
     Z100            :out std_logic;
     Z101            :out std_logic;
     Z102            :out std_logic;
     Z103            :out std_logic;
     Z104            :out std_logic;
     Z105            :out std_logic;
     Z106            :out std_logic;
     Z107            :out std_logic;
     Z108            :out std_logic;
     Z109            :out std_logic;
     Z110            :out std_logic;
     Z111            :out std_logic;
     Z112            :out std_logic;
     Z113            :out std_logic;
     Z114            :out std_logic;
     Z115            :out std_logic;
     Z116            :out std_logic;
     Z117            :out std_logic;
     Z118            :out std_logic;
     Z119            :out std_logic;
     Z120            :out std_logic;
     Z121            :out std_logic;
     Z122            :out std_logic;
     Z123            :out std_logic;
     Z124            :out std_logic;
     Z125            :out std_logic;
     Z126            :out std_logic;
     Z127            :out std_logic;
     Z128            :out std_logic;
     Z129            :out std_logic;
     Z130            :out std_logic;
     Z131            :out std_logic;
     Z132            :out std_logic;
     Z133            :out std_logic;
     Z134            :out std_logic;
     Z135            :out std_logic;
     Z136            :out std_logic;
     Z137            :out std_logic;
     Z138            :out std_logic;
     Z139            :out std_logic;
     Z140            :out std_logic;
     Z141            :out std_logic;
     Z142            :out std_logic;
     Z143            :out std_logic;
     Z144            :out std_logic;
     Z145            :out std_logic;
     Z146            :out std_logic;
     Z147            :out std_logic;
     Z148            :out std_logic;
     Z149            :out std_logic;
     Z150            :out std_logic;
     Z151            :out std_logic;
     Z152            :out std_logic;
     Z153            :out std_logic;
     Z154            :out std_logic;
     Z155            :out std_logic;
     Z156            :out std_logic;
     Z157            :out std_logic;
     Z158            :out std_logic;
     Z159            :out std_logic;
     Z160            :out std_logic;
     Z161            :out std_logic;
     Z162            :out std_logic;
     Z163            :out std_logic;
     Z164            :out std_logic;
     Z165            :out std_logic;
     Z166            :out std_logic;
     Z167            :out std_logic;
     Z168            :out std_logic;
     Z169            :out std_logic;
     Z170            :out std_logic;
     Z171            :out std_logic;
     Z172            :out std_logic;
     Z173            :out std_logic;
     Z174            :out std_logic;
     Z175            :out std_logic;
     Z176            :out std_logic;
     Z177            :out std_logic;
     Z178            :out std_logic;
     Z179            :out std_logic;
     Z180            :out std_logic;
     Z181            :out std_logic;
     Z182            :out std_logic;
     Z183            :out std_logic;
     Z184            :out std_logic;
     Z185            :out std_logic;
     Z186            :out std_logic;
     Z187            :out std_logic;
     Z188            :out std_logic;
     Z189            :out std_logic;
     Z190            :out std_logic;
     Z191            :out std_logic;
     Z192            :out std_logic;
     Z193            :out std_logic;
     Z194            :out std_logic;
     Z195            :out std_logic;
     Z196            :out std_logic;
     Z197            :out std_logic;
     Z198            :out std_logic;
     Z199            :out std_logic;
     Z200            :out std_logic;
     Z201            :out std_logic;
     Z202            :out std_logic;
     Z203            :out std_logic;
     Z204            :out std_logic;
     Z205            :out std_logic;
     Z206            :out std_logic;
     Z207            :out std_logic;
     Z208            :out std_logic;
     Z209            :out std_logic;
     Z210            :out std_logic;
     Z211            :out std_logic;
     Z212            :out std_logic;
     Z213            :out std_logic;
     Z214            :out std_logic;
     Z215            :out std_logic;
     Z216            :out std_logic;
     Z217            :out std_logic;
     Z218            :out std_logic;
     Z219            :out std_logic;
     Z220            :out std_logic;
     Z221            :out std_logic;
     Z222            :out std_logic;
     Z223            :out std_logic;
     Z224            :out std_logic;
     Z225            :out std_logic;
     Z226            :out std_logic;
     Z227            :out std_logic;
     Z228            :out std_logic;
     Z229            :out std_logic;
     Z230            :out std_logic;
     Z231            :out std_logic;
     Z232            :out std_logic;
     Z233            :out std_logic;
     Z234            :out std_logic;
     Z235            :out std_logic;
     Z236            :out std_logic;
     Z237            :out std_logic;
     Z238            :out std_logic;
     Z239            :out std_logic;
     Z240            :out std_logic;
     Z241            :out std_logic;
     Z242            :out std_logic;
     Z243            :out std_logic;
     Z244            :out std_logic;
     Z245            :out std_logic;
     Z246            :out std_logic;
     Z247            :out std_logic;
     Z248            :out std_logic;
     Z249            :out std_logic;
     Z250            :out std_logic;
     Z251            :out std_logic;
     Z252            :out std_logic;
     Z253            :out std_logic;
     Z254            :out std_logic;
     Z255            :out std_logic;
     Z256            :out std_logic;
     Z257            :out std_logic;
     Z258            :out std_logic;
     Z259            :out std_logic;
     Z260            :out std_logic;
     Z261            :out std_logic;
     Z262            :out std_logic;
     Z263            :out std_logic;
     Z264            :out std_logic;
     Z265            :out std_logic;
     Z266            :out std_logic;
     Z267            :out std_logic;
     Z268            :out std_logic;
     Z269            :out std_logic;
     Z270            :out std_logic;
     Z271            :out std_logic;
     Z272            :out std_logic;
     Z273            :out std_logic;
     Z274            :out std_logic;
     Z275            :out std_logic;
     Z276            :out std_logic;
     Z277            :out std_logic;
     Z278            :out std_logic;
     Z279            :out std_logic;
     Z280            :out std_logic;
     Z281            :out std_logic;
     Z282            :out std_logic;
     Z283            :out std_logic;
     Z284            :out std_logic;
     Z285            :out std_logic;
     Z286            :out std_logic;
     Z287            :out std_logic;
     Z288            :out std_logic;
     Z289            :out std_logic;
     Z290            :out std_logic;
     Z291            :out std_logic;
     Z292            :out std_logic;
     Z293            :out std_logic;
     Z294            :out std_logic;
     Z295            :out std_logic;
     Z296            :out std_logic;
     Z297            :out std_logic;
     Z298            :out std_logic;
     Z299            :out std_logic;
     Z300            :out std_logic;
     Z301            :out std_logic;
     Z302            :out std_logic;
     Z303            :out std_logic;
     Z304            :out std_logic;
     Z305            :out std_logic;
     Z306            :out std_logic;
     Z307            :out std_logic;
     Z308            :out std_logic;
     Z309            :out std_logic;
     Z310            :out std_logic;
     Z311            :out std_logic;
     Z312            :out std_logic;
     Z313            :out std_logic;
     Z314            :out std_logic;
     Z315            :out std_logic;
     Z316            :out std_logic;
     Z317            :out std_logic;
     Z318            :out std_logic;
     Z319            :out std_logic;
     Z320            :out std_logic;
     Z321            :out std_logic;
     Z322            :out std_logic;
     Z323            :out std_logic;
     Z324            :out std_logic;
     Z325            :out std_logic;
     Z326            :out std_logic;
     Z327            :out std_logic;
     Z328            :out std_logic;
     Z329            :out std_logic;
     Z330            :out std_logic;
     Z331            :out std_logic;
     Z332            :out std_logic;
     Z333            :out std_logic;
     Z334            :out std_logic;
     Z335            :out std_logic;
     Z336            :out std_logic;
     Z337            :out std_logic;
     Z338            :out std_logic;
     Z339            :out std_logic;
     Z340            :out std_logic;
     Z341            :out std_logic;
     Z342            :out std_logic;
     Z343            :out std_logic;
     Z344            :out std_logic;
     Z345            :out std_logic;
     Z346            :out std_logic;
     Z347            :out std_logic;
     Z348            :out std_logic;
     Z349            :out std_logic;
     Z350            :out std_logic;
     Z351            :out std_logic;
     Z352            :out std_logic;
     Z353            :out std_logic;
     Z354            :out std_logic;
     Z355            :out std_logic;
     Z356            :out std_logic;
     Z357            :out std_logic;
     Z358            :out std_logic;
     Z359            :out std_logic;
     Z360            :out std_logic;
     Z361            :out std_logic;
     Z362            :out std_logic;
     Z363            :out std_logic;
     Z364            :out std_logic;
     Z365            :out std_logic;
     Z366            :out std_logic;
     Z367            :out std_logic;
     Z368            :out std_logic;
     Z369            :out std_logic;
     Z370            :out std_logic;
     Z371            :out std_logic;
     Z372            :out std_logic;
     Z373            :out std_logic;
     Z374            :out std_logic;
     Z375            :out std_logic;
     Z376            :out std_logic;
     Z377            :out std_logic;
     Z378            :out std_logic;
     Z379            :out std_logic;
     Z380            :out std_logic;
     Z381            :out std_logic;
     Z382            :out std_logic;
     Z383            :out std_logic;
     Z384            :out std_logic;
     Z385            :out std_logic;
     Z386            :out std_logic;
     Z387            :out std_logic;
     Z388            :out std_logic;
     Z389            :out std_logic;
     Z390            :out std_logic;
     Z391            :out std_logic;
     Z392            :out std_logic;
     Z393            :out std_logic;
     Z394            :out std_logic;
     Z395            :out std_logic;
     Z396            :out std_logic;
     Z397            :out std_logic;
     Z398            :out std_logic;
     Z399            :out std_logic;
     Z400            :out std_logic;
     Z401            :out std_logic;
     Z402            :out std_logic;
     Z403            :out std_logic;
     Z404            :out std_logic;
     Z405            :out std_logic;
     Z406            :out std_logic;
     Z407            :out std_logic;
     Z408            :out std_logic;
     Z409            :out std_logic;
     Z410            :out std_logic;
     Z411            :out std_logic;
     Z412            :out std_logic;
     Z413            :out std_logic;
     Z414            :out std_logic;
     Z415            :out std_logic;
     Z416            :out std_logic;
     Z417            :out std_logic;
     Z418            :out std_logic;
     Z419            :out std_logic;
     Z420            :out std_logic;
     Z421            :out std_logic;
     Z422            :out std_logic;
     Z423            :out std_logic;
     Z424            :out std_logic;
     Z425            :out std_logic;
     Z426            :out std_logic;
     Z427            :out std_logic;
     Z428            :out std_logic;
     Z429            :out std_logic;
     Z430            :out std_logic;
     Z431            :out std_logic;
     Z432            :out std_logic;
     Z433            :out std_logic;
     Z434            :out std_logic;
     Z435            :out std_logic;
     Z436            :out std_logic;
     Z437            :out std_logic;
     Z438            :out std_logic;
     Z439            :out std_logic;
     Z440            :out std_logic;
     Z441            :out std_logic;
     Z442            :out std_logic;
     Z443            :out std_logic;
     Z444            :out std_logic;
     Z445            :out std_logic;
     Z446            :out std_logic;
     Z447            :out std_logic;
     Z448            :out std_logic;
     Z449            :out std_logic;
     Z450            :out std_logic;
     Z451            :out std_logic;
     Z452            :out std_logic;
     Z453            :out std_logic;
     Z454            :out std_logic;
     Z455            :out std_logic;
     Z456            :out std_logic;
     Z457            :out std_logic;
     Z458            :out std_logic;
     Z459            :out std_logic;
     Z460            :out std_logic;
     Z461            :out std_logic;
     Z462            :out std_logic;
     Z463            :out std_logic;
     Z464            :out std_logic;
     Z465            :out std_logic;
     Z466            :out std_logic;
     Z467            :out std_logic;
     Z468            :out std_logic;
     Z469            :out std_logic;
     Z470            :out std_logic;
     Z471            :out std_logic;
     Z472            :out std_logic;
     Z473            :out std_logic;
     Z474            :out std_logic;
     Z475            :out std_logic;
     Z476            :out std_logic;
     Z477            :out std_logic;
     Z478            :out std_logic;
     Z479            :out std_logic;
     Z480            :out std_logic;
     Z481            :out std_logic;
     Z482            :out std_logic;
     Z483            :out std_logic;
     Z484            :out std_logic;
     Z485            :out std_logic;
     Z486            :out std_logic;
     Z487            :out std_logic;
     Z488            :out std_logic;
     Z489            :out std_logic;
     Z490            :out std_logic;
     Z491            :out std_logic;
     Z492            :out std_logic;
     Z493            :out std_logic;
     Z494            :out std_logic;
     Z495            :out std_logic;
     Z496            :out std_logic;
     Z497            :out std_logic;
     Z498            :out std_logic;
     Z499            :out std_logic;
     Z500            :out std_logic;
     Z501            :out std_logic;
     Z502            :out std_logic;
     Z503            :out std_logic;
     Z504            :out std_logic;
     Z505            :out std_logic;
     Z506            :out std_logic;
     Z507            :out std_logic;
     Z508            :out std_logic;
     Z509            :out std_logic;
     Z510            :out std_logic;
     Z511            :out std_logic;
     Z512            :out std_logic;
     Z513            :out std_logic;
     Z514            :out std_logic;
     Z515            :out std_logic;
     Z516            :out std_logic;
     Z517            :out std_logic;
     Z518            :out std_logic;
     Z519            :out std_logic;
     Z520            :out std_logic;
     Z521            :out std_logic;
     Z522            :out std_logic;
     Z523            :out std_logic;
     Z524            :out std_logic;
     Z525            :out std_logic;
     Z526            :out std_logic;
     Z527            :out std_logic;
     Z528            :out std_logic;
     Z529            :out std_logic;
     Z530            :out std_logic;
     Z531            :out std_logic;
     Z532            :out std_logic;
     Z533            :out std_logic;
     Z534            :out std_logic;
     Z535            :out std_logic;
     Z536            :out std_logic;
     Z537            :out std_logic;
     Z538            :out std_logic;
     Z539            :out std_logic;
     Z540            :out std_logic;
     Z541            :out std_logic;
     Z542            :out std_logic;
     Z543            :out std_logic;
     Z544            :out std_logic;
     Z545            :out std_logic;
     Z546            :out std_logic;
     Z547            :out std_logic;
     Z548            :out std_logic;
     Z549            :out std_logic;
     Z550            :out std_logic;
     Z551            :out std_logic;
     Z552            :out std_logic;
     Z553            :out std_logic;
     Z554            :out std_logic;
     Z555            :out std_logic;
     Z556            :out std_logic;
     Z557            :out std_logic;
     Z558            :out std_logic;
     Z559            :out std_logic;
     Z560            :out std_logic;
     Z561            :out std_logic;
     Z562            :out std_logic;
     Z563            :out std_logic;
     Z564            :out std_logic;
     Z565            :out std_logic;
     Z566            :out std_logic;
     Z567            :out std_logic;
     Z568            :out std_logic;
     Z569            :out std_logic;
     Z570            :out std_logic;
     Z571            :out std_logic;
     Z572            :out std_logic;
     Z573            :out std_logic;
     Z574            :out std_logic;
     Z575            :out std_logic;
     Z576            :out std_logic;
     Z577            :out std_logic;
     Z578            :out std_logic;
     Z579            :out std_logic;
     Z580            :out std_logic;
     Z581            :out std_logic;
     Z582            :out std_logic;
     Z583            :out std_logic;
     Z584            :out std_logic;
     Z585            :out std_logic;
     Z586            :out std_logic;
     Z587            :out std_logic;
     Z588            :out std_logic;
     Z589            :out std_logic;
     Z590            :out std_logic;
     Z591            :out std_logic;
     Z592            :out std_logic;
     Z593            :out std_logic;
     Z594            :out std_logic;
     Z595            :out std_logic;
     Z596            :out std_logic;
     Z597            :out std_logic;
     Z598            :out std_logic;
     Z599            :out std_logic;
     Z600            :out std_logic;
     Z601            :out std_logic;
     Z602            :out std_logic;
     Z603            :out std_logic;
     Z604            :out std_logic;
     Z605            :out std_logic;
     Z606            :out std_logic;
     Z607            :out std_logic;
     Z608            :out std_logic;
     Z609            :out std_logic;
     Z610            :out std_logic;
     Z611            :out std_logic;
     Z612            :out std_logic;
     Z613            :out std_logic;
     Z614            :out std_logic;
     Z615            :out std_logic;
     Z616            :out std_logic;
     Z617            :out std_logic;
     Z618            :out std_logic;
     Z619            :out std_logic;
     Z620            :out std_logic;
     Z621            :out std_logic;
     Z622            :out std_logic;
     Z623            :out std_logic;
     Z624            :out std_logic;
     Z625            :out std_logic;
     Z626            :out std_logic;
     Z627            :out std_logic;
     Z628            :out std_logic;
     Z629            :out std_logic;
     Z630            :out std_logic;
     Z631            :out std_logic;
     Z632            :out std_logic;
     Z633            :out std_logic;
     Z634            :out std_logic;
     Z635            :out std_logic;
     Z636            :out std_logic;
     Z637            :out std_logic;
     Z638            :out std_logic;
     Z639            :out std_logic;
     Z640            :out std_logic;
     Z641            :out std_logic;
     Z642            :out std_logic;
     Z643            :out std_logic;
     Z644            :out std_logic;
     Z645            :out std_logic;
     Z646            :out std_logic;
     Z647            :out std_logic;
     Z648            :out std_logic;
     Z649            :out std_logic;
     Z650            :out std_logic;
     Z651            :out std_logic;
     Z652            :out std_logic;
     Z653            :out std_logic;
     Z654            :out std_logic;
     Z655            :out std_logic;
     Z656            :out std_logic;
     Z657            :out std_logic;
     Z658            :out std_logic;
     Z659            :out std_logic;
     Z660            :out std_logic;
     Z661            :out std_logic;
     Z662            :out std_logic;
     Z663            :out std_logic;
     Z664            :out std_logic;
     Z665            :out std_logic;
     Z666            :out std_logic;
     Z667            :out std_logic;
     Z668            :out std_logic;
     Z669            :out std_logic;
     Z670            :out std_logic;
     Z671            :out std_logic;
     Z672            :out std_logic;
     Z673            :out std_logic;
     Z674            :out std_logic;
     Z675            :out std_logic;
     Z676            :out std_logic;
     Z677            :out std_logic;
     Z678            :out std_logic;
     Z679            :out std_logic;
     Z680            :out std_logic;
     Z681            :out std_logic;
     Z682            :out std_logic;
     Z683            :out std_logic;
     Z684            :out std_logic;
     Z685            :out std_logic;
     Z686            :out std_logic;
     Z687            :out std_logic;
     Z688            :out std_logic;
     Z689            :out std_logic;
     Z690            :out std_logic;
     Z691            :out std_logic;
     Z692            :out std_logic;
     Z693            :out std_logic;
     Z694            :out std_logic;
     Z695            :out std_logic;
     Z696            :out std_logic;
     Z697            :out std_logic;
     Z698            :out std_logic;
     Z699            :out std_logic;
     Z700            :out std_logic;
     Z701            :out std_logic;
     Z702            :out std_logic;
     Z703            :out std_logic;
     Z704            :out std_logic;
     Z705            :out std_logic;
     Z706            :out std_logic;
     Z707            :out std_logic;
     Z708            :out std_logic;
     Z709            :out std_logic;
     Z710            :out std_logic;
     Z711            :out std_logic;
     Z712            :out std_logic;
     Z713            :out std_logic;
     Z714            :out std_logic;
     Z715            :out std_logic;
     Z716            :out std_logic;
     Z717            :out std_logic;
     Z718            :out std_logic;
     Z719            :out std_logic;
     Z720            :out std_logic;
     Z721            :out std_logic;
     Z722            :out std_logic;
     Z723            :out std_logic;
     Z724            :out std_logic;
     Z725            :out std_logic;
     Z726            :out std_logic;
     Z727            :out std_logic;
     Z728            :out std_logic;
     Z729            :out std_logic;
     Z730            :out std_logic;
     Z731            :out std_logic;
     Z732            :out std_logic;
     Z733            :out std_logic;
     Z734            :out std_logic;
     Z735            :out std_logic;
     Z736            :out std_logic;
     Z737            :out std_logic;
     Z738            :out std_logic;
     Z739            :out std_logic;
     Z740            :out std_logic;
     Z741            :out std_logic;
     Z742            :out std_logic;
     Z743            :out std_logic;
     Z744            :out std_logic;
     Z745            :out std_logic;
     Z746            :out std_logic;
     Z747            :out std_logic;
     Z748            :out std_logic;
     Z749            :out std_logic;
     Z750            :out std_logic;
     Z751            :out std_logic;
     Z752            :out std_logic;
     Z753            :out std_logic;
     Z754            :out std_logic;
     Z755            :out std_logic;
     Z756            :out std_logic;
     Z757            :out std_logic;
     Z758            :out std_logic;
     Z759            :out std_logic;
     Z760            :out std_logic;
     Z761            :out std_logic;
     Z762            :out std_logic;
     Z763            :out std_logic;
     Z764            :out std_logic;
     Z765            :out std_logic;
     Z766            :out std_logic;
     Z767            :out std_logic;
     Z768            :out std_logic;
     Z769            :out std_logic;
     Z770            :out std_logic;
     Z771            :out std_logic;
     Z772            :out std_logic;
     Z773            :out std_logic;
     Z774            :out std_logic;
     Z775            :out std_logic;
     Z776            :out std_logic;
     Z777            :out std_logic;
     Z778            :out std_logic;
     Z779            :out std_logic;
     Z780            :out std_logic;
     Z781            :out std_logic;
     Z782            :out std_logic;
     Z783            :out std_logic;
     Z784            :out std_logic;
     Z785            :out std_logic;
     Z786            :out std_logic;
     Z787            :out std_logic;
     Z788            :out std_logic;
     Z789            :out std_logic;
     Z790            :out std_logic;
     Z791            :out std_logic;
     Z792            :out std_logic;
     Z793            :out std_logic;
     Z794            :out std_logic;
     Z795            :out std_logic;
     Z796            :out std_logic;
     Z797            :out std_logic;
     Z798            :out std_logic;
     Z799            :out std_logic;
     Z800            :out std_logic;
     Z801            :out std_logic;
     Z802            :out std_logic;
     Z803            :out std_logic;
     Z804            :out std_logic;
     Z805            :out std_logic;
     Z806            :out std_logic;
     Z807            :out std_logic;
     Z808            :out std_logic;
     Z809            :out std_logic;
     Z810            :out std_logic;
     Z811            :out std_logic;
     Z812            :out std_logic;
     Z813            :out std_logic;
     Z814            :out std_logic;
     Z815            :out std_logic;
     Z816            :out std_logic;
     Z817            :out std_logic;
     Z818            :out std_logic;
     Z819            :out std_logic;
     Z820            :out std_logic;
     Z821            :out std_logic;
     Z822            :out std_logic;
     Z823            :out std_logic;
     Z824            :out std_logic;
     Z825            :out std_logic;
     Z826            :out std_logic;
     Z827            :out std_logic;
     Z828            :out std_logic;
     Z829            :out std_logic;
     Z830            :out std_logic;
     Z831            :out std_logic;
     Z832            :out std_logic;
     Z833            :out std_logic;
     Z834            :out std_logic;
     Z835            :out std_logic;
     Z836            :out std_logic;
     Z837            :out std_logic;
     Z838            :out std_logic;
     Z839            :out std_logic;
     Z840            :out std_logic;
     Z841            :out std_logic;
     Z842            :out std_logic;
     Z843            :out std_logic;
     Z844            :out std_logic;
     Z845            :out std_logic;
     Z846            :out std_logic;
     Z847            :out std_logic;
     Z848            :out std_logic;
     Z849            :out std_logic;
     Z850            :out std_logic;
     Z851            :out std_logic;
     Z852            :out std_logic;
     Z853            :out std_logic;
     Z854            :out std_logic;
     Z855            :out std_logic;
     Z856            :out std_logic;
     Z857            :out std_logic;
     Z858            :out std_logic;
     Z859            :out std_logic;
     Z860            :out std_logic;
     Z861            :out std_logic;
     Z862            :out std_logic;
     Z863            :out std_logic;
     Z864            :out std_logic;
     Z865            :out std_logic;
     Z866            :out std_logic;
     Z867            :out std_logic;
     Z868            :out std_logic;
     Z869            :out std_logic;
     Z870            :out std_logic;
     Z871            :out std_logic;
     Z872            :out std_logic;
     Z873            :out std_logic;
     Z874            :out std_logic;
     Z875            :out std_logic;
     Z876            :out std_logic;
     Z877            :out std_logic;
     Z878            :out std_logic;
     Z879            :out std_logic;
     Z880            :out std_logic;
     Z881            :out std_logic;
     Z882            :out std_logic;
     Z883            :out std_logic;
     Z884            :out std_logic;
     Z885            :out std_logic;
     Z886            :out std_logic;
     Z887            :out std_logic;
     Z888            :out std_logic;
     Z889            :out std_logic;
     Z890            :out std_logic;
     Z891            :out std_logic;
     Z892            :out std_logic;
     Z893            :out std_logic;
     Z894            :out std_logic;
     Z895            :out std_logic;
     Z896            :out std_logic;
     Z897            :out std_logic;
     Z898            :out std_logic;
     Z899            :out std_logic;
     Z900            :out std_logic;
     Z901            :out std_logic;
     Z902            :out std_logic;
     Z903            :out std_logic;
     Z904            :out std_logic;
     Z905            :out std_logic;
     Z906            :out std_logic;
     Z907            :out std_logic;
     Z908            :out std_logic;
     Z909            :out std_logic;
     Z910            :out std_logic;
     Z911            :out std_logic;
     Z912            :out std_logic;
     Z913            :out std_logic;
     Z914            :out std_logic;
     Z915            :out std_logic;
     Z916            :out std_logic;
     Z917            :out std_logic;
     Z918            :out std_logic;
     Z919            :out std_logic;
     Z920            :out std_logic;
     Z921            :out std_logic;
     Z922            :out std_logic;
     Z923            :out std_logic;
     Z924            :out std_logic;
     Z925            :out std_logic;
     Z926            :out std_logic;
     Z927            :out std_logic;
     Z928            :out std_logic;
     Z929            :out std_logic;
     Z930            :out std_logic;
     Z931            :out std_logic;
     Z932            :out std_logic;
     Z933            :out std_logic;
     Z934            :out std_logic;
     Z935            :out std_logic;
     Z936            :out std_logic;
     Z937            :out std_logic;
     Z938            :out std_logic;
     Z939            :out std_logic;
     Z940            :out std_logic;
     Z941            :out std_logic;
     Z942            :out std_logic;
     Z943            :out std_logic;
     Z944            :out std_logic;
     Z945            :out std_logic;
     Z946            :out std_logic;
     Z947            :out std_logic;
     Z948            :out std_logic;
     Z949            :out std_logic;
     Z950            :out std_logic;
     Z951            :out std_logic;
     Z952            :out std_logic;
     Z953            :out std_logic;
     Z954            :out std_logic;
     Z955            :out std_logic;
     Z956            :out std_logic;
     Z957            :out std_logic;
     Z958            :out std_logic;
     Z959            :out std_logic;
     Z960            :out std_logic;
     Z961            :out std_logic;
     Z962            :out std_logic;
     Z963            :out std_logic;
     Z964            :out std_logic;
     Z965            :out std_logic;
     Z966            :out std_logic;
     Z967            :out std_logic;
     Z968            :out std_logic;
     Z969            :out std_logic;
     Z970            :out std_logic;
     Z971            :out std_logic;
     Z972            :out std_logic;
     Z973            :out std_logic;
     Z974            :out std_logic;
     Z975            :out std_logic;
     Z976            :out std_logic;
     Z977            :out std_logic;
     Z978            :out std_logic;
     Z979            :out std_logic;
     Z980            :out std_logic;
     Z981            :out std_logic;
     Z982            :out std_logic;
     Z983            :out std_logic;
     Z984            :out std_logic;
     Z985            :out std_logic;
     Z986            :out std_logic;
     Z987            :out std_logic;
     Z988            :out std_logic;
     Z989            :out std_logic;
     Z990            :out std_logic;
     Z991            :out std_logic;
     Z992            :out std_logic;
     Z993            :out std_logic;
     Z994            :out std_logic;
     Z995            :out std_logic;
     Z996            :out std_logic;
     Z997            :out std_logic;
     Z998            :out std_logic;
     Z999            :out std_logic;
     Z1000            :out std_logic;
     Z1001            :out std_logic;
     Z1002            :out std_logic;
     Z1003            :out std_logic;
     Z1004            :out std_logic;
     Z1005            :out std_logic;
     Z1006            :out std_logic;
     Z1007            :out std_logic;
     Z1008            :out std_logic;
     Z1009            :out std_logic;
     Z1010            :out std_logic;
     Z1011            :out std_logic;
     Z1012            :out std_logic;
     Z1013            :out std_logic;
     Z1014            :out std_logic;
     Z1015            :out std_logic;
     Z1016            :out std_logic;
     Z1017            :out std_logic;
     Z1018            :out std_logic;
     Z1019            :out std_logic;
     Z1020            :out std_logic;
     Z1021            :out std_logic;
     Z1022            :out std_logic;
     Z1023            :out std_logic;
     Z1024            :out std_logic;
     Z1025            :out std_logic;
     Z1026            :out std_logic;
     Z1027            :out std_logic;
     Z1028            :out std_logic;
     Z1029            :out std_logic;
     Z1030            :out std_logic;
     Z1031            :out std_logic;
     Z1032            :out std_logic;
     Z1033            :out std_logic;
     Z1034            :out std_logic;
     Z1035            :out std_logic;
     Z1036            :out std_logic;
     Z1037            :out std_logic;
     Z1038            :out std_logic;
     Z1039            :out std_logic;
     Z1040            :out std_logic;
     Z1041            :out std_logic;
     Z1042            :out std_logic;
     Z1043            :out std_logic;
     Z1044            :out std_logic;
     Z1045            :out std_logic;
     Z1046            :out std_logic;
     Z1047            :out std_logic;
     Z1048            :out std_logic;
     Z1049            :out std_logic;
     Z1050            :out std_logic;
     Z1051            :out std_logic;
     Z1052            :out std_logic;
     Z1053            :out std_logic;
     Z1054            :out std_logic;
     Z1055            :out std_logic;
     Z1056            :out std_logic;
     Z1057            :out std_logic;
     Z1058            :out std_logic;
     Z1059            :out std_logic;
     Z1060            :out std_logic;
     Z1061            :out std_logic;
     Z1062            :out std_logic;
     Z1063            :out std_logic;
     Z1064            :out std_logic;
     Z1065            :out std_logic;
     Z1066            :out std_logic;
     Z1067            :out std_logic;
     Z1068            :out std_logic;
     Z1069            :out std_logic;
     Z1070            :out std_logic;
     Z1071            :out std_logic;
     Z1072            :out std_logic;
     Z1073            :out std_logic;
     Z1074            :out std_logic;
     Z1075            :out std_logic;
     Z1076            :out std_logic;
     Z1077            :out std_logic;
     Z1078            :out std_logic;
     Z1079            :out std_logic;
     Z1080            :out std_logic;
     Z1081            :out std_logic;
     Z1082            :out std_logic;
     Z1083            :out std_logic;
     Z1084            :out std_logic;
     Z1085            :out std_logic;
     Z1086            :out std_logic;
     Z1087            :out std_logic;
     Z1088            :out std_logic;
     Z1089            :out std_logic;
     Z1090            :out std_logic;
     Z1091            :out std_logic;
     Z1092            :out std_logic;
     Z1093            :out std_logic;
     Z1094            :out std_logic;
     Z1095            :out std_logic;
     Z1096            :out std_logic;
     Z1097            :out std_logic;
     Z1098            :out std_logic;
     Z1099            :out std_logic;
     Z1100            :out std_logic;
     Z1101            :out std_logic;
     Z1102            :out std_logic;
     Z1103            :out std_logic;
     Z1104            :out std_logic;
     Z1105            :out std_logic;
     Z1106            :out std_logic;
     Z1107            :out std_logic;
     Z1108            :out std_logic;
     Z1109            :out std_logic;
     Z1110            :out std_logic;
     Z1111            :out std_logic;
     Z1112            :out std_logic;
     Z1113            :out std_logic;
     Z1114            :out std_logic;
     Z1115            :out std_logic;
     Z1116            :out std_logic;
     Z1117            :out std_logic;
     Z1118            :out std_logic;
     Z1119            :out std_logic;
     Z1120            :out std_logic;
     Z1121            :out std_logic;
     Z1122            :out std_logic;
     Z1123            :out std_logic;
     Z1124            :out std_logic;
     Z1125            :out std_logic;
     Z1126            :out std_logic;
     Z1127            :out std_logic;
     Z1128            :out std_logic;
     Z1129            :out std_logic;
     Z1130            :out std_logic;
     Z1131            :out std_logic;
     Z1132            :out std_logic;
     Z1133            :out std_logic;
     Z1134            :out std_logic;
     Z1135            :out std_logic;
     Z1136            :out std_logic;
     Z1137            :out std_logic;
     Z1138            :out std_logic;
     Z1139            :out std_logic;
     Z1140            :out std_logic;
     Z1141            :out std_logic;
     Z1142            :out std_logic;
     Z1143            :out std_logic;
     Z1144            :out std_logic;
     Z1145            :out std_logic;
     Z1146            :out std_logic;
     Z1147            :out std_logic;
     Z1148            :out std_logic;
     Z1149            :out std_logic;
     Z1150            :out std_logic;
     Z1151            :out std_logic;
     Z1152            :out std_logic;
     Z1153            :out std_logic;
     Z1154            :out std_logic;
     Z1155            :out std_logic;
     Z1156            :out std_logic;
     Z1157            :out std_logic;
     Z1158            :out std_logic;
     Z1159            :out std_logic;
     Z1160            :out std_logic;
     Z1161            :out std_logic;
     Z1162            :out std_logic;
     Z1163            :out std_logic;
     Z1164            :out std_logic;
     Z1165            :out std_logic;
     Z1166            :out std_logic;
     Z1167            :out std_logic;
     Z1168            :out std_logic;
     Z1169            :out std_logic;
     Z1170            :out std_logic;
     Z1171            :out std_logic;
     Z1172            :out std_logic;
     Z1173            :out std_logic;
     Z1174            :out std_logic;
     Z1175            :out std_logic;
     Z1176            :out std_logic;
     Z1177            :out std_logic;
     Z1178            :out std_logic;
     Z1179            :out std_logic;
     Z1180            :out std_logic;
     Z1181            :out std_logic;
     Z1182            :out std_logic;
     Z1183            :out std_logic;
     Z1184            :out std_logic;
     Z1185            :out std_logic;
     Z1186            :out std_logic;
     Z1187            :out std_logic;
     Z1188            :out std_logic;
     Z1189            :out std_logic;
     Z1190            :out std_logic;
     Z1191            :out std_logic;
     Z1192            :out std_logic;
     Z1193            :out std_logic;
     Z1194            :out std_logic;
     Z1195            :out std_logic;
     Z1196            :out std_logic;
     Z1197            :out std_logic;
     Z1198            :out std_logic;
     Z1199            :out std_logic;
     Z1200            :out std_logic;
     Z1201            :out std_logic;
     Z1202            :out std_logic;
     Z1203            :out std_logic;
     Z1204            :out std_logic;
     Z1205            :out std_logic;
     Z1206            :out std_logic;
     Z1207            :out std_logic;
     Z1208            :out std_logic;
     Z1209            :out std_logic;
     Z1210            :out std_logic;
     Z1211            :out std_logic;
     Z1212            :out std_logic;
     Z1213            :out std_logic;
     Z1214            :out std_logic;
     Z1215            :out std_logic;
     Z1216            :out std_logic;
     Z1217            :out std_logic;
     Z1218            :out std_logic;
     Z1219            :out std_logic;
     Z1220            :out std_logic;
     Z1221            :out std_logic;
     Z1222            :out std_logic;
     Z1223            :out std_logic;
     Z1224            :out std_logic;
     Z1225            :out std_logic;
     Z1226            :out std_logic;
     Z1227            :out std_logic;
     Z1228            :out std_logic;
     Z1229            :out std_logic;
     Z1230            :out std_logic;
     Z1231            :out std_logic;
     Z1232            :out std_logic;
     Z1233            :out std_logic;
     Z1234            :out std_logic;
     Z1235            :out std_logic;
     Z1236            :out std_logic;
     Z1237            :out std_logic;
     Z1238            :out std_logic;
     Z1239            :out std_logic;
     Z1240            :out std_logic;
     Z1241            :out std_logic;
     Z1242            :out std_logic;
     Z1243            :out std_logic;
     Z1244            :out std_logic;
     Z1245            :out std_logic;
     Z1246            :out std_logic;
     Z1247            :out std_logic;
     Z1248            :out std_logic;
     Z1249            :out std_logic;
     Z1250            :out std_logic;
     Z1251            :out std_logic;
     Z1252            :out std_logic;
     Z1253            :out std_logic;
     Z1254            :out std_logic;
     Z1255            :out std_logic;
     Z1256            :out std_logic;
     Z1257            :out std_logic;
     Z1258            :out std_logic;
     Z1259            :out std_logic;
     Z1260            :out std_logic;
     Z1261            :out std_logic;
     Z1262            :out std_logic;
     Z1263            :out std_logic;
     Z1264            :out std_logic;
     Z1265            :out std_logic;
     Z1266            :out std_logic;
     Z1267            :out std_logic;
     Z1268            :out std_logic;
     Z1269            :out std_logic;
     Z1270            :out std_logic;
     Z1271            :out std_logic;
     Z1272            :out std_logic;
     Z1273            :out std_logic;
     Z1274            :out std_logic;
     Z1275            :out std_logic;
     Z1276            :out std_logic;
     Z1277            :out std_logic;
     Z1278            :out std_logic;
     Z1279            :out std_logic;
     Z1280            :out std_logic;
     Z1281            :out std_logic;
     Z1282            :out std_logic;
     Z1283            :out std_logic;
     Z1284            :out std_logic;
     Z1285            :out std_logic;
     Z1286            :out std_logic;
     Z1287            :out std_logic;
     Z1288            :out std_logic;
     Z1289            :out std_logic;
     Z1290            :out std_logic;
     Z1291            :out std_logic;
     Z1292            :out std_logic;
     Z1293            :out std_logic;
     Z1294            :out std_logic;
     Z1295            :out std_logic;
     Z1296            :out std_logic;
     Z1297            :out std_logic;
     Z1298            :out std_logic;
     Z1299            :out std_logic;
     Z1300            :out std_logic;
     Z1301            :out std_logic;
     Z1302            :out std_logic;
     Z1303            :out std_logic;
     Z1304            :out std_logic;
     Z1305            :out std_logic;
     Z1306            :out std_logic;
     Z1307            :out std_logic;
     Z1308            :out std_logic;
     Z1309            :out std_logic;
     Z1310            :out std_logic;
     Z1311            :out std_logic;
     Z1312            :out std_logic;
     Z1313            :out std_logic;
     Z1314            :out std_logic;
     Z1315            :out std_logic;
     Z1316            :out std_logic;
     Z1317            :out std_logic;
     Z1318            :out std_logic;
     Z1319            :out std_logic;
     Z1320            :out std_logic;
     Z1321            :out std_logic;
     Z1322            :out std_logic;
     Z1323            :out std_logic;
     Z1324            :out std_logic;
     Z1325            :out std_logic;
     Z1326            :out std_logic;
     Z1327            :out std_logic;
     Z1328            :out std_logic;
     Z1329            :out std_logic;
     Z1330            :out std_logic;
     Z1331            :out std_logic;
     Z1332            :out std_logic;
     Z1333            :out std_logic;
     Z1334            :out std_logic;
     Z1335            :out std_logic;
     Z1336            :out std_logic;
     Z1337            :out std_logic;
     Z1338            :out std_logic;
     Z1339            :out std_logic;
     Z1340            :out std_logic;
     Z1341            :out std_logic;
     Z1342            :out std_logic;
     Z1343            :out std_logic;
     Z1344            :out std_logic;
     Z1345            :out std_logic;
     Z1346            :out std_logic;
     Z1347            :out std_logic;
     Z1348            :out std_logic;
     Z1349            :out std_logic;
     Z1350            :out std_logic;
     Z1351            :out std_logic;
     Z1352            :out std_logic;
     Z1353            :out std_logic;
     Z1354            :out std_logic;
     Z1355            :out std_logic;
     Z1356            :out std_logic;
     Z1357            :out std_logic;
     Z1358            :out std_logic;
     Z1359            :out std_logic;
     Z1360            :out std_logic;
     Z1361            :out std_logic;
     Z1362            :out std_logic;
     Z1363            :out std_logic;
     Z1364            :out std_logic;
     Z1365            :out std_logic;
     Z1366            :out std_logic;
     Z1367            :out std_logic;
     Z1368            :out std_logic;
     Z1369            :out std_logic;
     Z1370            :out std_logic;
     Z1371            :out std_logic;
     Z1372            :out std_logic;
     Z1373            :out std_logic;
     Z1374            :out std_logic;
     Z1375            :out std_logic;
     Z1376            :out std_logic;
     Z1377            :out std_logic;
     Z1378            :out std_logic;
     Z1379            :out std_logic;
     Z1380            :out std_logic;
     Z1381            :out std_logic;
     Z1382            :out std_logic;
     Z1383            :out std_logic;
     Z1384            :out std_logic;
     Z1385            :out std_logic;
     Z1386            :out std_logic;
     Z1387            :out std_logic;
     Z1388            :out std_logic;
     Z1389            :out std_logic;
     Z1390            :out std_logic;
     Z1391            :out std_logic;
     Z1392            :out std_logic;
     Z1393            :out std_logic;
     Z1394            :out std_logic;
     Z1395            :out std_logic;
     Z1396            :out std_logic;
     Z1397            :out std_logic;
     Z1398            :out std_logic;
     Z1399            :out std_logic;
     Z1400            :out std_logic;
     Z1401            :out std_logic;
     Z1402            :out std_logic;
     Z1403            :out std_logic;
     Z1404            :out std_logic;
     Z1405            :out std_logic;
     Z1406            :out std_logic;
     Z1407            :out std_logic;
     Z1408            :out std_logic;
     Z1409            :out std_logic;
     Z1410            :out std_logic;
     Z1411            :out std_logic;
     Z1412            :out std_logic;
     Z1413            :out std_logic;
     Z1414            :out std_logic;
     Z1415            :out std_logic;
     Z1416            :out std_logic;
     Z1417            :out std_logic;
     Z1418            :out std_logic;
     Z1419            :out std_logic;
     Z1420            :out std_logic;
     Z1421            :out std_logic;
     Z1422            :out std_logic;
     Z1423            :out std_logic;
     Z1424            :out std_logic;
     Z1425            :out std_logic;
     Z1426            :out std_logic;
     Z1427            :out std_logic;
     Z1428            :out std_logic;
     Z1429            :out std_logic;
     Z1430            :out std_logic;
     Z1431            :out std_logic;
     Z1432            :out std_logic;
     Z1433            :out std_logic;
     Z1434            :out std_logic;
     Z1435            :out std_logic;
     Z1436            :out std_logic;
     Z1437            :out std_logic;
     Z1438            :out std_logic;
     Z1439            :out std_logic;
     Z1440            :out std_logic;
     Z1441            :out std_logic;
     Z1442            :out std_logic;
     Z1443            :out std_logic;
     Z1444            :out std_logic;
     Z1445            :out std_logic;
     Z1446            :out std_logic;
     Z1447            :out std_logic;
     Z1448            :out std_logic;
     Z1449            :out std_logic;
     Z1450            :out std_logic;
     Z1451            :out std_logic;
     Z1452            :out std_logic;
     Z1453            :out std_logic;
     Z1454            :out std_logic;
     Z1455            :out std_logic;
     Z1456            :out std_logic;
     Z1457            :out std_logic;
     Z1458            :out std_logic;
     Z1459            :out std_logic;
     Z1460            :out std_logic;
     Z1461            :out std_logic;
     Z1462            :out std_logic;
     Z1463            :out std_logic;
     Z1464            :out std_logic;
     Z1465            :out std_logic;
     Z1466            :out std_logic;
     Z1467            :out std_logic;
     Z1468            :out std_logic;
     Z1469            :out std_logic;
     Z1470            :out std_logic;
     Z1471            :out std_logic;
     Z1472            :out std_logic;
     Z1473            :out std_logic;
     Z1474            :out std_logic;
     Z1475            :out std_logic;
     Z1476            :out std_logic;
     Z1477            :out std_logic;
     Z1478            :out std_logic;
     Z1479            :out std_logic;
     Z1480            :out std_logic;
     Z1481            :out std_logic;
     Z1482            :out std_logic;
     Z1483            :out std_logic;
     Z1484            :out std_logic;
     Z1485            :out std_logic;
     Z1486            :out std_logic;
     Z1487            :out std_logic;
     Z1488            :out std_logic;
     Z1489            :out std_logic;
     Z1490            :out std_logic;
     Z1491            :out std_logic;
     Z1492            :out std_logic;
     Z1493            :out std_logic;
     Z1494            :out std_logic;
     Z1495            :out std_logic;
     Z1496            :out std_logic;
     Z1497            :out std_logic;
     Z1498            :out std_logic;
     Z1499            :out std_logic;
     Z1500            :out std_logic;
     Z1501            :out std_logic;
     Z1502            :out std_logic;
     Z1503            :out std_logic;
     Z1504            :out std_logic;
     Z1505            :out std_logic;
     Z1506            :out std_logic;
     Z1507            :out std_logic;
     Z1508            :out std_logic;
     Z1509            :out std_logic;
     Z1510            :out std_logic;
     Z1511            :out std_logic;
     Z1512            :out std_logic;
     Z1513            :out std_logic;
     Z1514            :out std_logic;
     Z1515            :out std_logic;
     Z1516            :out std_logic;
     Z1517            :out std_logic;
     Z1518            :out std_logic;
     Z1519            :out std_logic;
     Z1520            :out std_logic;
     Z1521            :out std_logic;
     Z1522            :out std_logic;
     Z1523            :out std_logic;
     Z1524            :out std_logic;
     Z1525            :out std_logic;
     Z1526            :out std_logic;
     Z1527            :out std_logic;
     Z1528            :out std_logic;
     Z1529            :out std_logic;
     Z1530            :out std_logic;
     Z1531            :out std_logic;
     Z1532            :out std_logic;
     Z1533            :out std_logic;
     Z1534            :out std_logic;
     Z1535            :out std_logic;
     Z1536            :out std_logic;
     Z1537            :out std_logic;
     Z1538            :out std_logic;
     Z1539            :out std_logic;
     Z1540            :out std_logic;
     Z1541            :out std_logic;
     Z1542            :out std_logic;
     Z1543            :out std_logic;
     Z1544            :out std_logic;
     Z1545            :out std_logic;
     Z1546            :out std_logic;
     Z1547            :out std_logic;
     Z1548            :out std_logic;
     Z1549            :out std_logic;
     Z1550            :out std_logic;
     Z1551            :out std_logic;
     Z1552            :out std_logic;
     Z1553            :out std_logic;
     Z1554            :out std_logic;
     Z1555            :out std_logic;
     Z1556            :out std_logic;
     Z1557            :out std_logic;
     Z1558            :out std_logic;
     Z1559            :out std_logic;
     Z1560            :out std_logic;
     Z1561            :out std_logic;
     Z1562            :out std_logic;
     Z1563            :out std_logic;
     Z1564            :out std_logic;
     Z1565            :out std_logic;
     Z1566            :out std_logic;
     Z1567            :out std_logic;
     Z1568            :out std_logic;
     Z1569            :out std_logic;
     Z1570            :out std_logic;
     Z1571            :out std_logic;
     Z1572            :out std_logic;
     Z1573            :out std_logic;
     Z1574            :out std_logic;
     Z1575            :out std_logic;
     Z1576            :out std_logic;
     Z1577            :out std_logic;
     Z1578            :out std_logic;
     Z1579            :out std_logic;
     Z1580            :out std_logic;
     Z1581            :out std_logic;
     Z1582            :out std_logic;
     Z1583            :out std_logic;
     Z1584            :out std_logic;
     Z1585            :out std_logic;
     Z1586            :out std_logic;
     Z1587            :out std_logic;
     Z1588            :out std_logic;
     Z1589            :out std_logic;
     Z1590            :out std_logic;
     Z1591            :out std_logic;
     Z1592            :out std_logic;
     Z1593            :out std_logic;
     Z1594            :out std_logic;
     Z1595            :out std_logic;
     Z1596            :out std_logic;
     Z1597            :out std_logic;
     Z1598            :out std_logic;
     Z1599            :out std_logic;
     Z1600            :out std_logic;
     Z1601            :out std_logic;
     Z1602            :out std_logic;
     Z1603            :out std_logic;
     Z1604            :out std_logic;
     Z1605            :out std_logic;
     Z1606            :out std_logic;
     Z1607            :out std_logic;
     Z1608            :out std_logic;
     Z1609            :out std_logic;
     Z1610            :out std_logic;
     Z1611            :out std_logic;
     Z1612            :out std_logic;
     Z1613            :out std_logic;
     Z1614            :out std_logic;
     Z1615            :out std_logic;
     Z1616            :out std_logic;
     Z1617            :out std_logic;
     Z1618            :out std_logic;
     Z1619            :out std_logic;
     Z1620            :out std_logic;
     Z1621            :out std_logic;
     Z1622            :out std_logic;
     Z1623            :out std_logic;
     Z1624            :out std_logic;
     Z1625            :out std_logic;
     Z1626            :out std_logic;
     Z1627            :out std_logic;
     Z1628            :out std_logic;
     Z1629            :out std_logic;
     Z1630            :out std_logic;
     Z1631            :out std_logic;
     Z1632            :out std_logic;
     Z1633            :out std_logic;
     Z1634            :out std_logic;
     Z1635            :out std_logic;
     Z1636            :out std_logic;
     Z1637            :out std_logic;
     Z1638            :out std_logic;
     Z1639            :out std_logic;
     Z1640            :out std_logic;
     Z1641            :out std_logic;
     Z1642            :out std_logic;
     Z1643            :out std_logic;
     Z1644            :out std_logic;
     Z1645            :out std_logic;
     Z1646            :out std_logic;
     Z1647            :out std_logic;
     Z1648            :out std_logic;
     Z1649            :out std_logic;
     Z1650            :out std_logic;
     Z1651            :out std_logic;
     Z1652            :out std_logic;
     Z1653            :out std_logic;
     Z1654            :out std_logic;
     Z1655            :out std_logic;
     Z1656            :out std_logic;
     Z1657            :out std_logic;
     Z1658            :out std_logic;
     Z1659            :out std_logic;
     Z1660            :out std_logic;
     Z1661            :out std_logic;
     Z1662            :out std_logic;
     Z1663            :out std_logic;
     Z1664            :out std_logic;
     Z1665            :out std_logic;
     Z1666            :out std_logic;
     Z1667            :out std_logic;
     Z1668            :out std_logic;
     Z1669            :out std_logic;
     Z1670            :out std_logic;
     Z1671            :out std_logic;
     Z1672            :out std_logic;
     Z1673            :out std_logic;
     Z1674            :out std_logic;
     Z1675            :out std_logic;
     Z1676            :out std_logic;
     Z1677            :out std_logic;
     Z1678            :out std_logic;
     Z1679            :out std_logic;
     Z1680            :out std_logic;
     Z1681            :out std_logic;
     Z1682            :out std_logic;
     Z1683            :out std_logic;
     Z1684            :out std_logic;
     Z1685            :out std_logic;
     Z1686            :out std_logic;
     Z1687            :out std_logic;
     Z1688            :out std_logic;
     Z1689            :out std_logic;
     Z1690            :out std_logic;
     Z1691            :out std_logic;
     Z1692            :out std_logic;
     Z1693            :out std_logic;
     Z1694            :out std_logic;
     Z1695            :out std_logic;
     Z1696            :out std_logic;
     Z1697            :out std_logic;
     Z1698            :out std_logic;
     Z1699            :out std_logic;
     Z1700            :out std_logic;
     Z1701            :out std_logic;
     Z1702            :out std_logic;
     Z1703            :out std_logic;
     Z1704            :out std_logic;
     Z1705            :out std_logic;
     Z1706            :out std_logic;
     Z1707            :out std_logic;
     Z1708            :out std_logic;
     Z1709            :out std_logic;
     Z1710            :out std_logic;
     Z1711            :out std_logic;
     Z1712            :out std_logic;
     Z1713            :out std_logic;
     Z1714            :out std_logic;
     Z1715            :out std_logic;
     Z1716            :out std_logic;
     Z1717            :out std_logic;
     Z1718            :out std_logic;
     Z1719            :out std_logic;
     Z1720            :out std_logic;
     Z1721            :out std_logic;
     Z1722            :out std_logic;
     Z1723            :out std_logic;
     Z1724            :out std_logic;
     Z1725            :out std_logic;
     Z1726            :out std_logic;
     Z1727            :out std_logic;
     Z1728            :out std_logic;
     Z1729            :out std_logic;
     Z1730            :out std_logic;
     Z1731            :out std_logic;
     Z1732            :out std_logic;
     Z1733            :out std_logic;
     Z1734            :out std_logic;
     Z1735            :out std_logic;
     Z1736            :out std_logic;
     Z1737            :out std_logic;
     Z1738            :out std_logic;
     Z1739            :out std_logic;
     Z1740            :out std_logic;
     Z1741            :out std_logic;
     Z1742            :out std_logic;
     Z1743            :out std_logic;
     Z1744            :out std_logic;
     Z1745            :out std_logic;
     Z1746            :out std_logic;
     Z1747            :out std_logic;
     Z1748            :out std_logic;
     Z1749            :out std_logic;
     Z1750            :out std_logic;
     Z1751            :out std_logic;
     Z1752            :out std_logic;
     Z1753            :out std_logic;
     Z1754            :out std_logic;
     Z1755            :out std_logic;
     Z1756            :out std_logic;
     Z1757            :out std_logic;
     Z1758            :out std_logic;
     Z1759            :out std_logic;
     Z1760            :out std_logic;
     Z1761            :out std_logic;
     Z1762            :out std_logic;
     Z1763            :out std_logic;
     Z1764            :out std_logic;
     Z1765            :out std_logic;
     Z1766            :out std_logic;
     Z1767            :out std_logic;
     Z1768            :out std_logic;
     Z1769            :out std_logic;
     Z1770            :out std_logic;
     Z1771            :out std_logic;
     Z1772            :out std_logic;
     Z1773            :out std_logic;
     Z1774            :out std_logic;
     Z1775            :out std_logic;
     Z1776            :out std_logic;
     Z1777            :out std_logic;
     Z1778            :out std_logic;
     Z1779            :out std_logic;
     Z1780            :out std_logic;
     Z1781            :out std_logic;
     Z1782            :out std_logic;
     Z1783            :out std_logic;
     Z1784            :out std_logic;
     Z1785            :out std_logic;
     Z1786            :out std_logic;
     Z1787            :out std_logic;
     Z1788            :out std_logic;
     Z1789            :out std_logic;
     Z1790            :out std_logic;
     Z1791            :out std_logic;
     Z1792            :out std_logic;
     Z1793            :out std_logic;
     Z1794            :out std_logic;
     Z1795            :out std_logic;
     Z1796            :out std_logic;
     Z1797            :out std_logic;
     Z1798            :out std_logic;
     Z1799            :out std_logic;
     Z1800            :out std_logic;
     Z1801            :out std_logic;
     Z1802            :out std_logic;
     Z1803            :out std_logic;
     Z1804            :out std_logic;
     Z1805            :out std_logic;
     Z1806            :out std_logic;
     Z1807            :out std_logic;
     Z1808            :out std_logic;
     Z1809            :out std_logic;
     Z1810            :out std_logic;
     Z1811            :out std_logic;
     Z1812            :out std_logic;
     Z1813            :out std_logic;
     Z1814            :out std_logic;
     Z1815            :out std_logic;
     Z1816            :out std_logic;
     Z1817            :out std_logic;
     Z1818            :out std_logic;
     Z1819            :out std_logic;
     Z1820            :out std_logic;
     Z1821            :out std_logic;
     Z1822            :out std_logic;
     Z1823            :out std_logic;
     Z1824            :out std_logic;
     Z1825            :out std_logic;
     Z1826            :out std_logic;
     Z1827            :out std_logic;
     Z1828            :out std_logic;
     Z1829            :out std_logic;
     Z1830            :out std_logic;
     Z1831            :out std_logic;
     Z1832            :out std_logic;
     Z1833            :out std_logic;
     Z1834            :out std_logic;
     Z1835            :out std_logic;
     Z1836            :out std_logic;
     Z1837            :out std_logic;
     Z1838            :out std_logic;
     Z1839            :out std_logic;
     Z1840            :out std_logic;
     Z1841            :out std_logic;
     Z1842            :out std_logic;
     Z1843            :out std_logic;
     Z1844            :out std_logic;
     Z1845            :out std_logic;
     Z1846            :out std_logic;
     Z1847            :out std_logic;
     Z1848            :out std_logic;
     Z1849            :out std_logic;
     Z1850            :out std_logic;
     Z1851            :out std_logic;
     Z1852            :out std_logic;
     Z1853            :out std_logic;
     Z1854            :out std_logic;
     Z1855            :out std_logic;
     Z1856            :out std_logic;
     Z1857            :out std_logic;
     Z1858            :out std_logic;
     Z1859            :out std_logic;
     Z1860            :out std_logic;
     Z1861            :out std_logic;
     Z1862            :out std_logic;
     Z1863            :out std_logic;
     Z1864            :out std_logic;
     Z1865            :out std_logic;
     Z1866            :out std_logic;
     Z1867            :out std_logic;
     Z1868            :out std_logic;
     Z1869            :out std_logic;
     Z1870            :out std_logic;
     Z1871            :out std_logic;
     Z1872            :out std_logic;
     Z1873            :out std_logic;
     Z1874            :out std_logic;
     Z1875            :out std_logic;
     Z1876            :out std_logic;
     Z1877            :out std_logic;
     Z1878            :out std_logic;
     Z1879            :out std_logic;
     Z1880            :out std_logic;
     Z1881            :out std_logic;
     Z1882            :out std_logic;
     Z1883            :out std_logic;
     Z1884            :out std_logic;
     Z1885            :out std_logic;
     Z1886            :out std_logic;
     Z1887            :out std_logic;
     Z1888            :out std_logic;
     Z1889            :out std_logic;
     Z1890            :out std_logic;
     Z1891            :out std_logic;
     Z1892            :out std_logic;
     Z1893            :out std_logic;
     Z1894            :out std_logic;
     Z1895            :out std_logic;
     Z1896            :out std_logic;
     Z1897            :out std_logic;
     Z1898            :out std_logic;
     Z1899            :out std_logic;
     Z1900            :out std_logic;
     Z1901            :out std_logic;
     Z1902            :out std_logic;
     Z1903            :out std_logic;
     Z1904            :out std_logic;
     Z1905            :out std_logic;
     Z1906            :out std_logic;
     Z1907            :out std_logic;
     Z1908            :out std_logic;
     Z1909            :out std_logic;
     Z1910            :out std_logic;
     Z1911            :out std_logic;
     Z1912            :out std_logic;
     Z1913            :out std_logic;
     Z1914            :out std_logic;
     Z1915            :out std_logic;
     Z1916            :out std_logic;
     Z1917            :out std_logic;
     Z1918            :out std_logic;
     Z1919            :out std_logic;
     Z1920            :out std_logic;
     Z1921            :out std_logic;
     Z1922            :out std_logic;
     Z1923            :out std_logic;
     Z1924            :out std_logic;
     Z1925            :out std_logic;
     Z1926            :out std_logic;
     Z1927            :out std_logic;
     Z1928            :out std_logic;
     Z1929            :out std_logic;
     Z1930            :out std_logic;
     Z1931            :out std_logic;
     Z1932            :out std_logic;
     Z1933            :out std_logic;
     Z1934            :out std_logic;
     Z1935            :out std_logic;
     Z1936            :out std_logic;
     Z1937            :out std_logic;
     Z1938            :out std_logic;
     Z1939            :out std_logic;
     Z1940            :out std_logic;
     Z1941            :out std_logic;
     Z1942            :out std_logic;
     Z1943            :out std_logic;
     Z1944            :out std_logic;
     Z1945            :out std_logic;
     Z1946            :out std_logic;
     Z1947            :out std_logic;
     Z1948            :out std_logic;
     Z1949            :out std_logic;
     Z1950            :out std_logic;
     Z1951            :out std_logic;
     Z1952            :out std_logic;
     Z1953            :out std_logic;
     Z1954            :out std_logic;
     Z1955            :out std_logic;
     Z1956            :out std_logic;
     Z1957            :out std_logic;
     Z1958            :out std_logic;
     Z1959            :out std_logic;
     Z1960            :out std_logic;
     Z1961            :out std_logic;
     Z1962            :out std_logic;
     Z1963            :out std_logic;
     Z1964            :out std_logic;
     Z1965            :out std_logic;
     Z1966            :out std_logic;
     Z1967            :out std_logic;
     Z1968            :out std_logic;
     Z1969            :out std_logic;
     Z1970            :out std_logic;
     Z1971            :out std_logic;
     Z1972            :out std_logic;
     Z1973            :out std_logic;
     Z1974            :out std_logic;
     Z1975            :out std_logic;
     Z1976            :out std_logic;
     Z1977            :out std_logic;
     Z1978            :out std_logic;
     Z1979            :out std_logic;
     Z1980            :out std_logic;
     Z1981            :out std_logic;
     Z1982            :out std_logic;
     Z1983            :out std_logic;
     Z1984            :out std_logic;
     Z1985            :out std_logic;
     Z1986            :out std_logic;
     Z1987            :out std_logic;
     Z1988            :out std_logic;
     Z1989            :out std_logic;
     Z1990            :out std_logic;
     Z1991            :out std_logic;
     Z1992            :out std_logic;
     Z1993            :out std_logic;
     Z1994            :out std_logic;
     Z1995            :out std_logic;
     Z1996            :out std_logic;
     Z1997            :out std_logic;
     Z1998            :out std_logic;
     Z1999            :out std_logic;
     Z2000            :out std_logic;
     Z2001            :out std_logic;
     Z2002            :out std_logic;
     Z2003            :out std_logic;
     Z2004            :out std_logic;
     Z2005            :out std_logic;
     Z2006            :out std_logic;
     Z2007            :out std_logic;
     Z2008            :out std_logic;
     Z2009            :out std_logic;
     Z2010            :out std_logic;
     Z2011            :out std_logic;
     Z2012            :out std_logic;
     Z2013            :out std_logic;
     Z2014            :out std_logic;
     Z2015            :out std_logic;
     Z2016            :out std_logic;
     Z2017            :out std_logic;
     Z2018            :out std_logic;
     Z2019            :out std_logic;
     Z2020            :out std_logic;
     Z2021            :out std_logic;
     Z2022            :out std_logic;
     Z2023            :out std_logic;
     Z2024            :out std_logic;
     Z2025            :out std_logic;
     Z2026            :out std_logic;
     Z2027            :out std_logic;
     Z2028            :out std_logic;
     Z2029            :out std_logic;
     Z2030            :out std_logic;
     Z2031            :out std_logic;
     Z2032            :out std_logic;
     Z2033            :out std_logic;
     Z2034            :out std_logic;
     Z2035            :out std_logic;
     Z2036            :out std_logic;
     Z2037            :out std_logic;
     Z2038            :out std_logic;
     Z2039            :out std_logic;
     Z2040            :out std_logic;
     Z2041            :out std_logic;
     Z2042            :out std_logic;
     Z2043            :out std_logic;
     Z2044            :out std_logic;
     Z2045            :out std_logic;
     Z2046            :out std_logic;
     Z2047            :out std_logic;
     Z2048            :out std_logic;
     Z2049            :out std_logic;
     Z2050            :out std_logic;
     Z2051            :out std_logic;
     Z2052            :out std_logic;
     Z2053            :out std_logic;
     Z2054            :out std_logic;
     Z2055            :out std_logic;
     Z2056            :out std_logic;
     Z2057            :out std_logic;
     Z2058            :out std_logic;
     Z2059            :out std_logic;
     Z2060            :out std_logic;
     Z2061            :out std_logic;
     Z2062            :out std_logic;
     Z2063            :out std_logic;
     Z2064            :out std_logic;
     Z2065            :out std_logic;
     Z2066            :out std_logic;
     Z2067            :out std_logic;
     Z2068            :out std_logic;
     Z2069            :out std_logic;
     Z2070            :out std_logic;
     Z2071            :out std_logic;
     Z2072            :out std_logic;
     Z2073            :out std_logic;
     Z2074            :out std_logic;
     Z2075            :out std_logic;
     Z2076            :out std_logic;
     Z2077            :out std_logic;
     Z2078            :out std_logic;
     Z2079            :out std_logic;
     Z2080            :out std_logic;
     Z2081            :out std_logic;
     Z2082            :out std_logic;
     Z2083            :out std_logic;
     Z2084            :out std_logic;
     Z2085            :out std_logic;
     Z2086            :out std_logic;
     Z2087            :out std_logic;
     Z2088            :out std_logic;
     Z2089            :out std_logic;
     Z2090            :out std_logic;
     Z2091            :out std_logic;
     Z2092            :out std_logic;
     Z2093            :out std_logic;
     Z2094            :out std_logic;
     Z2095            :out std_logic;
     Z2096            :out std_logic;
     Z2097            :out std_logic;
     Z2098            :out std_logic;
     Z2099            :out std_logic;
     Z2100            :out std_logic;
     Z2101            :out std_logic;
     Z2102            :out std_logic;
     Z2103            :out std_logic;
     Z2104            :out std_logic;
     Z2105            :out std_logic;
     Z2106            :out std_logic;
     Z2107            :out std_logic;
     Z2108            :out std_logic;
     Z2109            :out std_logic;
     Z2110            :out std_logic;
     Z2111            :out std_logic;
     Z2112            :out std_logic;
     Z2113            :out std_logic;
     Z2114            :out std_logic;
     Z2115            :out std_logic;
     Z2116            :out std_logic;
     Z2117            :out std_logic;
     Z2118            :out std_logic;
     Z2119            :out std_logic;
     Z2120            :out std_logic;
     Z2121            :out std_logic;
     Z2122            :out std_logic;
     Z2123            :out std_logic;
     Z2124            :out std_logic;
     Z2125            :out std_logic;
     Z2126            :out std_logic;
     Z2127            :out std_logic;
     Z2128            :out std_logic;
     Z2129            :out std_logic;
     Z2130            :out std_logic;
     Z2131            :out std_logic;
     Z2132            :out std_logic;
     Z2133            :out std_logic;
     Z2134            :out std_logic;
     Z2135            :out std_logic;
     Z2136            :out std_logic;
     Z2137            :out std_logic;
     Z2138            :out std_logic;
     Z2139            :out std_logic;
     Z2140            :out std_logic;
     Z2141            :out std_logic;
     Z2142            :out std_logic;
     Z2143            :out std_logic;
     Z2144            :out std_logic;
     Z2145            :out std_logic;
     Z2146            :out std_logic;
     Z2147            :out std_logic;
     Z2148            :out std_logic;
     Z2149            :out std_logic;
     Z2150            :out std_logic;
     Z2151            :out std_logic;
     Z2152            :out std_logic;
     Z2153            :out std_logic;
     Z2154            :out std_logic;
     Z2155            :out std_logic;
     Z2156            :out std_logic;
     Z2157            :out std_logic;
     Z2158            :out std_logic;
     Z2159            :out std_logic;
     Z2160            :out std_logic;
     Z2161            :out std_logic;
     Z2162            :out std_logic;
     Z2163            :out std_logic;
     Z2164            :out std_logic;
     Z2165            :out std_logic;
     Z2166            :out std_logic;
     Z2167            :out std_logic;
     Z2168            :out std_logic;
     Z2169            :out std_logic;
     Z2170            :out std_logic;
     Z2171            :out std_logic;
     Z2172            :out std_logic;
     Z2173            :out std_logic;
     Z2174            :out std_logic;
     Z2175            :out std_logic;
     Z2176            :out std_logic;
     Z2177            :out std_logic;
     Z2178            :out std_logic;
     Z2179            :out std_logic;
     Z2180            :out std_logic;
     Z2181            :out std_logic;
     Z2182            :out std_logic;
     Z2183            :out std_logic;
     Z2184            :out std_logic;
     Z2185            :out std_logic;
     Z2186            :out std_logic;
     Z2187            :out std_logic;
     Z2188            :out std_logic;
     Z2189            :out std_logic;
     Z2190            :out std_logic;
     Z2191            :out std_logic;
     Z2192            :out std_logic;
     Z2193            :out std_logic;
     Z2194            :out std_logic;
     Z2195            :out std_logic;
     Z2196            :out std_logic;
     Z2197            :out std_logic;
     Z2198            :out std_logic;
     Z2199            :out std_logic;
     Z2200            :out std_logic;
     Z2201            :out std_logic;
     Z2202            :out std_logic;
     Z2203            :out std_logic;
     Z2204            :out std_logic;
     Z2205            :out std_logic;
     Z2206            :out std_logic;
     Z2207            :out std_logic;
     Z2208            :out std_logic;
     Z2209            :out std_logic;
     Z2210            :out std_logic;
     Z2211            :out std_logic;
     Z2212            :out std_logic;
     Z2213            :out std_logic;
     Z2214            :out std_logic;
     Z2215            :out std_logic;
     Z2216            :out std_logic;
     Z2217            :out std_logic;
     Z2218            :out std_logic;
     Z2219            :out std_logic;
     Z2220            :out std_logic;
     Z2221            :out std_logic;
     Z2222            :out std_logic;
     Z2223            :out std_logic;
     Z2224            :out std_logic;
     Z2225            :out std_logic;
     Z2226            :out std_logic;
     Z2227            :out std_logic;
     Z2228            :out std_logic;
     Z2229            :out std_logic;
     Z2230            :out std_logic;
     Z2231            :out std_logic;
     Z2232            :out std_logic;
     Z2233            :out std_logic;
     Z2234            :out std_logic;
     Z2235            :out std_logic;
     Z2236            :out std_logic;
     Z2237            :out std_logic;
     Z2238            :out std_logic;
     Z2239            :out std_logic;
     Z2240            :out std_logic;
     Z2241            :out std_logic;
     Z2242            :out std_logic;
     Z2243            :out std_logic;
     Z2244            :out std_logic;
     Z2245            :out std_logic;
     Z2246            :out std_logic;
     Z2247            :out std_logic;
     Z2248            :out std_logic;
     Z2249            :out std_logic;
     Z2250            :out std_logic;
     Z2251            :out std_logic;
     Z2252            :out std_logic;
     Z2253            :out std_logic;
     Z2254            :out std_logic;
     Z2255            :out std_logic;
     Z2256            :out std_logic;
     Z2257            :out std_logic;
     Z2258            :out std_logic;
     Z2259            :out std_logic;
     Z2260            :out std_logic;
     Z2261            :out std_logic;
     Z2262            :out std_logic;
     Z2263            :out std_logic;
     Z2264            :out std_logic;
     Z2265            :out std_logic;
     Z2266            :out std_logic;
     Z2267            :out std_logic;
     Z2268            :out std_logic;
     Z2269            :out std_logic;
     Z2270            :out std_logic;
     Z2271            :out std_logic;
     Z2272            :out std_logic;
     Z2273            :out std_logic;
     Z2274            :out std_logic;
     Z2275            :out std_logic;
     Z2276            :out std_logic;
     Z2277            :out std_logic;
     Z2278            :out std_logic;
     Z2279            :out std_logic;
     Z2280            :out std_logic;
     Z2281            :out std_logic;
     Z2282            :out std_logic;
     Z2283            :out std_logic;
     Z2284            :out std_logic;
     Z2285            :out std_logic;
     Z2286            :out std_logic;
     Z2287            :out std_logic;
     Z2288            :out std_logic;
     Z2289            :out std_logic;
     Z2290            :out std_logic;
     Z2291            :out std_logic;
     Z2292            :out std_logic;
     Z2293            :out std_logic;
     Z2294            :out std_logic;
     Z2295            :out std_logic;
     Z2296            :out std_logic;
     Z2297            :out std_logic;
     Z2298            :out std_logic;
     Z2299            :out std_logic;
     Z2300            :out std_logic;
     Z2301            :out std_logic;
     Z2302            :out std_logic;
     Z2303            :out std_logic;
     Z2304            :out std_logic;
     num_iter         :out std_logic_vector(4 downto 0);
     end_decoder      :out std_logic
);
END;
ARCHITECTURE decoder_arch OF decoder IS

----------------------------- Declaration des components -------------------
 COMPONENT ldpc is PORT(
     clk,rst,start_vn,start_cn   :in std_logic;
     Lc1              :in std_logic_vector(8 DOWNTO 0);
     Lc2              :in std_logic_vector(8 DOWNTO 0);
     Lc3              :in std_logic_vector(8 DOWNTO 0);
     Lc4              :in std_logic_vector(8 DOWNTO 0);
     Lc5              :in std_logic_vector(8 DOWNTO 0);
     Lc6              :in std_logic_vector(8 DOWNTO 0);
     Lc7              :in std_logic_vector(8 DOWNTO 0);
     Lc8              :in std_logic_vector(8 DOWNTO 0);
     Lc9              :in std_logic_vector(8 DOWNTO 0);
     Lc10              :in std_logic_vector(8 DOWNTO 0);
     Lc11              :in std_logic_vector(8 DOWNTO 0);
     Lc12              :in std_logic_vector(8 DOWNTO 0);
     Lc13              :in std_logic_vector(8 DOWNTO 0);
     Lc14              :in std_logic_vector(8 DOWNTO 0);
     Lc15              :in std_logic_vector(8 DOWNTO 0);
     Lc16              :in std_logic_vector(8 DOWNTO 0);
     Lc17              :in std_logic_vector(8 DOWNTO 0);
     Lc18              :in std_logic_vector(8 DOWNTO 0);
     Lc19              :in std_logic_vector(8 DOWNTO 0);
     Lc20              :in std_logic_vector(8 DOWNTO 0);
     Lc21              :in std_logic_vector(8 DOWNTO 0);
     Lc22              :in std_logic_vector(8 DOWNTO 0);
     Lc23              :in std_logic_vector(8 DOWNTO 0);
     Lc24              :in std_logic_vector(8 DOWNTO 0);
     Lc25              :in std_logic_vector(8 DOWNTO 0);
     Lc26              :in std_logic_vector(8 DOWNTO 0);
     Lc27              :in std_logic_vector(8 DOWNTO 0);
     Lc28              :in std_logic_vector(8 DOWNTO 0);
     Lc29              :in std_logic_vector(8 DOWNTO 0);
     Lc30              :in std_logic_vector(8 DOWNTO 0);
     Lc31              :in std_logic_vector(8 DOWNTO 0);
     Lc32              :in std_logic_vector(8 DOWNTO 0);
     Lc33              :in std_logic_vector(8 DOWNTO 0);
     Lc34              :in std_logic_vector(8 DOWNTO 0);
     Lc35              :in std_logic_vector(8 DOWNTO 0);
     Lc36              :in std_logic_vector(8 DOWNTO 0);
     Lc37              :in std_logic_vector(8 DOWNTO 0);
     Lc38              :in std_logic_vector(8 DOWNTO 0);
     Lc39              :in std_logic_vector(8 DOWNTO 0);
     Lc40              :in std_logic_vector(8 DOWNTO 0);
     Lc41              :in std_logic_vector(8 DOWNTO 0);
     Lc42              :in std_logic_vector(8 DOWNTO 0);
     Lc43              :in std_logic_vector(8 DOWNTO 0);
     Lc44              :in std_logic_vector(8 DOWNTO 0);
     Lc45              :in std_logic_vector(8 DOWNTO 0);
     Lc46              :in std_logic_vector(8 DOWNTO 0);
     Lc47              :in std_logic_vector(8 DOWNTO 0);
     Lc48              :in std_logic_vector(8 DOWNTO 0);
     Lc49              :in std_logic_vector(8 DOWNTO 0);
     Lc50              :in std_logic_vector(8 DOWNTO 0);
     Lc51              :in std_logic_vector(8 DOWNTO 0);
     Lc52              :in std_logic_vector(8 DOWNTO 0);
     Lc53              :in std_logic_vector(8 DOWNTO 0);
     Lc54              :in std_logic_vector(8 DOWNTO 0);
     Lc55              :in std_logic_vector(8 DOWNTO 0);
     Lc56              :in std_logic_vector(8 DOWNTO 0);
     Lc57              :in std_logic_vector(8 DOWNTO 0);
     Lc58              :in std_logic_vector(8 DOWNTO 0);
     Lc59              :in std_logic_vector(8 DOWNTO 0);
     Lc60              :in std_logic_vector(8 DOWNTO 0);
     Lc61              :in std_logic_vector(8 DOWNTO 0);
     Lc62              :in std_logic_vector(8 DOWNTO 0);
     Lc63              :in std_logic_vector(8 DOWNTO 0);
     Lc64              :in std_logic_vector(8 DOWNTO 0);
     Lc65              :in std_logic_vector(8 DOWNTO 0);
     Lc66              :in std_logic_vector(8 DOWNTO 0);
     Lc67              :in std_logic_vector(8 DOWNTO 0);
     Lc68              :in std_logic_vector(8 DOWNTO 0);
     Lc69              :in std_logic_vector(8 DOWNTO 0);
     Lc70              :in std_logic_vector(8 DOWNTO 0);
     Lc71              :in std_logic_vector(8 DOWNTO 0);
     Lc72              :in std_logic_vector(8 DOWNTO 0);
     Lc73              :in std_logic_vector(8 DOWNTO 0);
     Lc74              :in std_logic_vector(8 DOWNTO 0);
     Lc75              :in std_logic_vector(8 DOWNTO 0);
     Lc76              :in std_logic_vector(8 DOWNTO 0);
     Lc77              :in std_logic_vector(8 DOWNTO 0);
     Lc78              :in std_logic_vector(8 DOWNTO 0);
     Lc79              :in std_logic_vector(8 DOWNTO 0);
     Lc80              :in std_logic_vector(8 DOWNTO 0);
     Lc81              :in std_logic_vector(8 DOWNTO 0);
     Lc82              :in std_logic_vector(8 DOWNTO 0);
     Lc83              :in std_logic_vector(8 DOWNTO 0);
     Lc84              :in std_logic_vector(8 DOWNTO 0);
     Lc85              :in std_logic_vector(8 DOWNTO 0);
     Lc86              :in std_logic_vector(8 DOWNTO 0);
     Lc87              :in std_logic_vector(8 DOWNTO 0);
     Lc88              :in std_logic_vector(8 DOWNTO 0);
     Lc89              :in std_logic_vector(8 DOWNTO 0);
     Lc90              :in std_logic_vector(8 DOWNTO 0);
     Lc91              :in std_logic_vector(8 DOWNTO 0);
     Lc92              :in std_logic_vector(8 DOWNTO 0);
     Lc93              :in std_logic_vector(8 DOWNTO 0);
     Lc94              :in std_logic_vector(8 DOWNTO 0);
     Lc95              :in std_logic_vector(8 DOWNTO 0);
     Lc96              :in std_logic_vector(8 DOWNTO 0);
     Lc97              :in std_logic_vector(8 DOWNTO 0);
     Lc98              :in std_logic_vector(8 DOWNTO 0);
     Lc99              :in std_logic_vector(8 DOWNTO 0);
     Lc100              :in std_logic_vector(8 DOWNTO 0);
     Lc101              :in std_logic_vector(8 DOWNTO 0);
     Lc102              :in std_logic_vector(8 DOWNTO 0);
     Lc103              :in std_logic_vector(8 DOWNTO 0);
     Lc104              :in std_logic_vector(8 DOWNTO 0);
     Lc105              :in std_logic_vector(8 DOWNTO 0);
     Lc106              :in std_logic_vector(8 DOWNTO 0);
     Lc107              :in std_logic_vector(8 DOWNTO 0);
     Lc108              :in std_logic_vector(8 DOWNTO 0);
     Lc109              :in std_logic_vector(8 DOWNTO 0);
     Lc110              :in std_logic_vector(8 DOWNTO 0);
     Lc111              :in std_logic_vector(8 DOWNTO 0);
     Lc112              :in std_logic_vector(8 DOWNTO 0);
     Lc113              :in std_logic_vector(8 DOWNTO 0);
     Lc114              :in std_logic_vector(8 DOWNTO 0);
     Lc115              :in std_logic_vector(8 DOWNTO 0);
     Lc116              :in std_logic_vector(8 DOWNTO 0);
     Lc117              :in std_logic_vector(8 DOWNTO 0);
     Lc118              :in std_logic_vector(8 DOWNTO 0);
     Lc119              :in std_logic_vector(8 DOWNTO 0);
     Lc120              :in std_logic_vector(8 DOWNTO 0);
     Lc121              :in std_logic_vector(8 DOWNTO 0);
     Lc122              :in std_logic_vector(8 DOWNTO 0);
     Lc123              :in std_logic_vector(8 DOWNTO 0);
     Lc124              :in std_logic_vector(8 DOWNTO 0);
     Lc125              :in std_logic_vector(8 DOWNTO 0);
     Lc126              :in std_logic_vector(8 DOWNTO 0);
     Lc127              :in std_logic_vector(8 DOWNTO 0);
     Lc128              :in std_logic_vector(8 DOWNTO 0);
     Lc129              :in std_logic_vector(8 DOWNTO 0);
     Lc130              :in std_logic_vector(8 DOWNTO 0);
     Lc131              :in std_logic_vector(8 DOWNTO 0);
     Lc132              :in std_logic_vector(8 DOWNTO 0);
     Lc133              :in std_logic_vector(8 DOWNTO 0);
     Lc134              :in std_logic_vector(8 DOWNTO 0);
     Lc135              :in std_logic_vector(8 DOWNTO 0);
     Lc136              :in std_logic_vector(8 DOWNTO 0);
     Lc137              :in std_logic_vector(8 DOWNTO 0);
     Lc138              :in std_logic_vector(8 DOWNTO 0);
     Lc139              :in std_logic_vector(8 DOWNTO 0);
     Lc140              :in std_logic_vector(8 DOWNTO 0);
     Lc141              :in std_logic_vector(8 DOWNTO 0);
     Lc142              :in std_logic_vector(8 DOWNTO 0);
     Lc143              :in std_logic_vector(8 DOWNTO 0);
     Lc144              :in std_logic_vector(8 DOWNTO 0);
     Lc145              :in std_logic_vector(8 DOWNTO 0);
     Lc146              :in std_logic_vector(8 DOWNTO 0);
     Lc147              :in std_logic_vector(8 DOWNTO 0);
     Lc148              :in std_logic_vector(8 DOWNTO 0);
     Lc149              :in std_logic_vector(8 DOWNTO 0);
     Lc150              :in std_logic_vector(8 DOWNTO 0);
     Lc151              :in std_logic_vector(8 DOWNTO 0);
     Lc152              :in std_logic_vector(8 DOWNTO 0);
     Lc153              :in std_logic_vector(8 DOWNTO 0);
     Lc154              :in std_logic_vector(8 DOWNTO 0);
     Lc155              :in std_logic_vector(8 DOWNTO 0);
     Lc156              :in std_logic_vector(8 DOWNTO 0);
     Lc157              :in std_logic_vector(8 DOWNTO 0);
     Lc158              :in std_logic_vector(8 DOWNTO 0);
     Lc159              :in std_logic_vector(8 DOWNTO 0);
     Lc160              :in std_logic_vector(8 DOWNTO 0);
     Lc161              :in std_logic_vector(8 DOWNTO 0);
     Lc162              :in std_logic_vector(8 DOWNTO 0);
     Lc163              :in std_logic_vector(8 DOWNTO 0);
     Lc164              :in std_logic_vector(8 DOWNTO 0);
     Lc165              :in std_logic_vector(8 DOWNTO 0);
     Lc166              :in std_logic_vector(8 DOWNTO 0);
     Lc167              :in std_logic_vector(8 DOWNTO 0);
     Lc168              :in std_logic_vector(8 DOWNTO 0);
     Lc169              :in std_logic_vector(8 DOWNTO 0);
     Lc170              :in std_logic_vector(8 DOWNTO 0);
     Lc171              :in std_logic_vector(8 DOWNTO 0);
     Lc172              :in std_logic_vector(8 DOWNTO 0);
     Lc173              :in std_logic_vector(8 DOWNTO 0);
     Lc174              :in std_logic_vector(8 DOWNTO 0);
     Lc175              :in std_logic_vector(8 DOWNTO 0);
     Lc176              :in std_logic_vector(8 DOWNTO 0);
     Lc177              :in std_logic_vector(8 DOWNTO 0);
     Lc178              :in std_logic_vector(8 DOWNTO 0);
     Lc179              :in std_logic_vector(8 DOWNTO 0);
     Lc180              :in std_logic_vector(8 DOWNTO 0);
     Lc181              :in std_logic_vector(8 DOWNTO 0);
     Lc182              :in std_logic_vector(8 DOWNTO 0);
     Lc183              :in std_logic_vector(8 DOWNTO 0);
     Lc184              :in std_logic_vector(8 DOWNTO 0);
     Lc185              :in std_logic_vector(8 DOWNTO 0);
     Lc186              :in std_logic_vector(8 DOWNTO 0);
     Lc187              :in std_logic_vector(8 DOWNTO 0);
     Lc188              :in std_logic_vector(8 DOWNTO 0);
     Lc189              :in std_logic_vector(8 DOWNTO 0);
     Lc190              :in std_logic_vector(8 DOWNTO 0);
     Lc191              :in std_logic_vector(8 DOWNTO 0);
     Lc192              :in std_logic_vector(8 DOWNTO 0);
     Lc193              :in std_logic_vector(8 DOWNTO 0);
     Lc194              :in std_logic_vector(8 DOWNTO 0);
     Lc195              :in std_logic_vector(8 DOWNTO 0);
     Lc196              :in std_logic_vector(8 DOWNTO 0);
     Lc197              :in std_logic_vector(8 DOWNTO 0);
     Lc198              :in std_logic_vector(8 DOWNTO 0);
     Lc199              :in std_logic_vector(8 DOWNTO 0);
     Lc200              :in std_logic_vector(8 DOWNTO 0);
     Lc201              :in std_logic_vector(8 DOWNTO 0);
     Lc202              :in std_logic_vector(8 DOWNTO 0);
     Lc203              :in std_logic_vector(8 DOWNTO 0);
     Lc204              :in std_logic_vector(8 DOWNTO 0);
     Lc205              :in std_logic_vector(8 DOWNTO 0);
     Lc206              :in std_logic_vector(8 DOWNTO 0);
     Lc207              :in std_logic_vector(8 DOWNTO 0);
     Lc208              :in std_logic_vector(8 DOWNTO 0);
     Lc209              :in std_logic_vector(8 DOWNTO 0);
     Lc210              :in std_logic_vector(8 DOWNTO 0);
     Lc211              :in std_logic_vector(8 DOWNTO 0);
     Lc212              :in std_logic_vector(8 DOWNTO 0);
     Lc213              :in std_logic_vector(8 DOWNTO 0);
     Lc214              :in std_logic_vector(8 DOWNTO 0);
     Lc215              :in std_logic_vector(8 DOWNTO 0);
     Lc216              :in std_logic_vector(8 DOWNTO 0);
     Lc217              :in std_logic_vector(8 DOWNTO 0);
     Lc218              :in std_logic_vector(8 DOWNTO 0);
     Lc219              :in std_logic_vector(8 DOWNTO 0);
     Lc220              :in std_logic_vector(8 DOWNTO 0);
     Lc221              :in std_logic_vector(8 DOWNTO 0);
     Lc222              :in std_logic_vector(8 DOWNTO 0);
     Lc223              :in std_logic_vector(8 DOWNTO 0);
     Lc224              :in std_logic_vector(8 DOWNTO 0);
     Lc225              :in std_logic_vector(8 DOWNTO 0);
     Lc226              :in std_logic_vector(8 DOWNTO 0);
     Lc227              :in std_logic_vector(8 DOWNTO 0);
     Lc228              :in std_logic_vector(8 DOWNTO 0);
     Lc229              :in std_logic_vector(8 DOWNTO 0);
     Lc230              :in std_logic_vector(8 DOWNTO 0);
     Lc231              :in std_logic_vector(8 DOWNTO 0);
     Lc232              :in std_logic_vector(8 DOWNTO 0);
     Lc233              :in std_logic_vector(8 DOWNTO 0);
     Lc234              :in std_logic_vector(8 DOWNTO 0);
     Lc235              :in std_logic_vector(8 DOWNTO 0);
     Lc236              :in std_logic_vector(8 DOWNTO 0);
     Lc237              :in std_logic_vector(8 DOWNTO 0);
     Lc238              :in std_logic_vector(8 DOWNTO 0);
     Lc239              :in std_logic_vector(8 DOWNTO 0);
     Lc240              :in std_logic_vector(8 DOWNTO 0);
     Lc241              :in std_logic_vector(8 DOWNTO 0);
     Lc242              :in std_logic_vector(8 DOWNTO 0);
     Lc243              :in std_logic_vector(8 DOWNTO 0);
     Lc244              :in std_logic_vector(8 DOWNTO 0);
     Lc245              :in std_logic_vector(8 DOWNTO 0);
     Lc246              :in std_logic_vector(8 DOWNTO 0);
     Lc247              :in std_logic_vector(8 DOWNTO 0);
     Lc248              :in std_logic_vector(8 DOWNTO 0);
     Lc249              :in std_logic_vector(8 DOWNTO 0);
     Lc250              :in std_logic_vector(8 DOWNTO 0);
     Lc251              :in std_logic_vector(8 DOWNTO 0);
     Lc252              :in std_logic_vector(8 DOWNTO 0);
     Lc253              :in std_logic_vector(8 DOWNTO 0);
     Lc254              :in std_logic_vector(8 DOWNTO 0);
     Lc255              :in std_logic_vector(8 DOWNTO 0);
     Lc256              :in std_logic_vector(8 DOWNTO 0);
     Lc257              :in std_logic_vector(8 DOWNTO 0);
     Lc258              :in std_logic_vector(8 DOWNTO 0);
     Lc259              :in std_logic_vector(8 DOWNTO 0);
     Lc260              :in std_logic_vector(8 DOWNTO 0);
     Lc261              :in std_logic_vector(8 DOWNTO 0);
     Lc262              :in std_logic_vector(8 DOWNTO 0);
     Lc263              :in std_logic_vector(8 DOWNTO 0);
     Lc264              :in std_logic_vector(8 DOWNTO 0);
     Lc265              :in std_logic_vector(8 DOWNTO 0);
     Lc266              :in std_logic_vector(8 DOWNTO 0);
     Lc267              :in std_logic_vector(8 DOWNTO 0);
     Lc268              :in std_logic_vector(8 DOWNTO 0);
     Lc269              :in std_logic_vector(8 DOWNTO 0);
     Lc270              :in std_logic_vector(8 DOWNTO 0);
     Lc271              :in std_logic_vector(8 DOWNTO 0);
     Lc272              :in std_logic_vector(8 DOWNTO 0);
     Lc273              :in std_logic_vector(8 DOWNTO 0);
     Lc274              :in std_logic_vector(8 DOWNTO 0);
     Lc275              :in std_logic_vector(8 DOWNTO 0);
     Lc276              :in std_logic_vector(8 DOWNTO 0);
     Lc277              :in std_logic_vector(8 DOWNTO 0);
     Lc278              :in std_logic_vector(8 DOWNTO 0);
     Lc279              :in std_logic_vector(8 DOWNTO 0);
     Lc280              :in std_logic_vector(8 DOWNTO 0);
     Lc281              :in std_logic_vector(8 DOWNTO 0);
     Lc282              :in std_logic_vector(8 DOWNTO 0);
     Lc283              :in std_logic_vector(8 DOWNTO 0);
     Lc284              :in std_logic_vector(8 DOWNTO 0);
     Lc285              :in std_logic_vector(8 DOWNTO 0);
     Lc286              :in std_logic_vector(8 DOWNTO 0);
     Lc287              :in std_logic_vector(8 DOWNTO 0);
     Lc288              :in std_logic_vector(8 DOWNTO 0);
     Lc289              :in std_logic_vector(8 DOWNTO 0);
     Lc290              :in std_logic_vector(8 DOWNTO 0);
     Lc291              :in std_logic_vector(8 DOWNTO 0);
     Lc292              :in std_logic_vector(8 DOWNTO 0);
     Lc293              :in std_logic_vector(8 DOWNTO 0);
     Lc294              :in std_logic_vector(8 DOWNTO 0);
     Lc295              :in std_logic_vector(8 DOWNTO 0);
     Lc296              :in std_logic_vector(8 DOWNTO 0);
     Lc297              :in std_logic_vector(8 DOWNTO 0);
     Lc298              :in std_logic_vector(8 DOWNTO 0);
     Lc299              :in std_logic_vector(8 DOWNTO 0);
     Lc300              :in std_logic_vector(8 DOWNTO 0);
     Lc301              :in std_logic_vector(8 DOWNTO 0);
     Lc302              :in std_logic_vector(8 DOWNTO 0);
     Lc303              :in std_logic_vector(8 DOWNTO 0);
     Lc304              :in std_logic_vector(8 DOWNTO 0);
     Lc305              :in std_logic_vector(8 DOWNTO 0);
     Lc306              :in std_logic_vector(8 DOWNTO 0);
     Lc307              :in std_logic_vector(8 DOWNTO 0);
     Lc308              :in std_logic_vector(8 DOWNTO 0);
     Lc309              :in std_logic_vector(8 DOWNTO 0);
     Lc310              :in std_logic_vector(8 DOWNTO 0);
     Lc311              :in std_logic_vector(8 DOWNTO 0);
     Lc312              :in std_logic_vector(8 DOWNTO 0);
     Lc313              :in std_logic_vector(8 DOWNTO 0);
     Lc314              :in std_logic_vector(8 DOWNTO 0);
     Lc315              :in std_logic_vector(8 DOWNTO 0);
     Lc316              :in std_logic_vector(8 DOWNTO 0);
     Lc317              :in std_logic_vector(8 DOWNTO 0);
     Lc318              :in std_logic_vector(8 DOWNTO 0);
     Lc319              :in std_logic_vector(8 DOWNTO 0);
     Lc320              :in std_logic_vector(8 DOWNTO 0);
     Lc321              :in std_logic_vector(8 DOWNTO 0);
     Lc322              :in std_logic_vector(8 DOWNTO 0);
     Lc323              :in std_logic_vector(8 DOWNTO 0);
     Lc324              :in std_logic_vector(8 DOWNTO 0);
     Lc325              :in std_logic_vector(8 DOWNTO 0);
     Lc326              :in std_logic_vector(8 DOWNTO 0);
     Lc327              :in std_logic_vector(8 DOWNTO 0);
     Lc328              :in std_logic_vector(8 DOWNTO 0);
     Lc329              :in std_logic_vector(8 DOWNTO 0);
     Lc330              :in std_logic_vector(8 DOWNTO 0);
     Lc331              :in std_logic_vector(8 DOWNTO 0);
     Lc332              :in std_logic_vector(8 DOWNTO 0);
     Lc333              :in std_logic_vector(8 DOWNTO 0);
     Lc334              :in std_logic_vector(8 DOWNTO 0);
     Lc335              :in std_logic_vector(8 DOWNTO 0);
     Lc336              :in std_logic_vector(8 DOWNTO 0);
     Lc337              :in std_logic_vector(8 DOWNTO 0);
     Lc338              :in std_logic_vector(8 DOWNTO 0);
     Lc339              :in std_logic_vector(8 DOWNTO 0);
     Lc340              :in std_logic_vector(8 DOWNTO 0);
     Lc341              :in std_logic_vector(8 DOWNTO 0);
     Lc342              :in std_logic_vector(8 DOWNTO 0);
     Lc343              :in std_logic_vector(8 DOWNTO 0);
     Lc344              :in std_logic_vector(8 DOWNTO 0);
     Lc345              :in std_logic_vector(8 DOWNTO 0);
     Lc346              :in std_logic_vector(8 DOWNTO 0);
     Lc347              :in std_logic_vector(8 DOWNTO 0);
     Lc348              :in std_logic_vector(8 DOWNTO 0);
     Lc349              :in std_logic_vector(8 DOWNTO 0);
     Lc350              :in std_logic_vector(8 DOWNTO 0);
     Lc351              :in std_logic_vector(8 DOWNTO 0);
     Lc352              :in std_logic_vector(8 DOWNTO 0);
     Lc353              :in std_logic_vector(8 DOWNTO 0);
     Lc354              :in std_logic_vector(8 DOWNTO 0);
     Lc355              :in std_logic_vector(8 DOWNTO 0);
     Lc356              :in std_logic_vector(8 DOWNTO 0);
     Lc357              :in std_logic_vector(8 DOWNTO 0);
     Lc358              :in std_logic_vector(8 DOWNTO 0);
     Lc359              :in std_logic_vector(8 DOWNTO 0);
     Lc360              :in std_logic_vector(8 DOWNTO 0);
     Lc361              :in std_logic_vector(8 DOWNTO 0);
     Lc362              :in std_logic_vector(8 DOWNTO 0);
     Lc363              :in std_logic_vector(8 DOWNTO 0);
     Lc364              :in std_logic_vector(8 DOWNTO 0);
     Lc365              :in std_logic_vector(8 DOWNTO 0);
     Lc366              :in std_logic_vector(8 DOWNTO 0);
     Lc367              :in std_logic_vector(8 DOWNTO 0);
     Lc368              :in std_logic_vector(8 DOWNTO 0);
     Lc369              :in std_logic_vector(8 DOWNTO 0);
     Lc370              :in std_logic_vector(8 DOWNTO 0);
     Lc371              :in std_logic_vector(8 DOWNTO 0);
     Lc372              :in std_logic_vector(8 DOWNTO 0);
     Lc373              :in std_logic_vector(8 DOWNTO 0);
     Lc374              :in std_logic_vector(8 DOWNTO 0);
     Lc375              :in std_logic_vector(8 DOWNTO 0);
     Lc376              :in std_logic_vector(8 DOWNTO 0);
     Lc377              :in std_logic_vector(8 DOWNTO 0);
     Lc378              :in std_logic_vector(8 DOWNTO 0);
     Lc379              :in std_logic_vector(8 DOWNTO 0);
     Lc380              :in std_logic_vector(8 DOWNTO 0);
     Lc381              :in std_logic_vector(8 DOWNTO 0);
     Lc382              :in std_logic_vector(8 DOWNTO 0);
     Lc383              :in std_logic_vector(8 DOWNTO 0);
     Lc384              :in std_logic_vector(8 DOWNTO 0);
     Lc385              :in std_logic_vector(8 DOWNTO 0);
     Lc386              :in std_logic_vector(8 DOWNTO 0);
     Lc387              :in std_logic_vector(8 DOWNTO 0);
     Lc388              :in std_logic_vector(8 DOWNTO 0);
     Lc389              :in std_logic_vector(8 DOWNTO 0);
     Lc390              :in std_logic_vector(8 DOWNTO 0);
     Lc391              :in std_logic_vector(8 DOWNTO 0);
     Lc392              :in std_logic_vector(8 DOWNTO 0);
     Lc393              :in std_logic_vector(8 DOWNTO 0);
     Lc394              :in std_logic_vector(8 DOWNTO 0);
     Lc395              :in std_logic_vector(8 DOWNTO 0);
     Lc396              :in std_logic_vector(8 DOWNTO 0);
     Lc397              :in std_logic_vector(8 DOWNTO 0);
     Lc398              :in std_logic_vector(8 DOWNTO 0);
     Lc399              :in std_logic_vector(8 DOWNTO 0);
     Lc400              :in std_logic_vector(8 DOWNTO 0);
     Lc401              :in std_logic_vector(8 DOWNTO 0);
     Lc402              :in std_logic_vector(8 DOWNTO 0);
     Lc403              :in std_logic_vector(8 DOWNTO 0);
     Lc404              :in std_logic_vector(8 DOWNTO 0);
     Lc405              :in std_logic_vector(8 DOWNTO 0);
     Lc406              :in std_logic_vector(8 DOWNTO 0);
     Lc407              :in std_logic_vector(8 DOWNTO 0);
     Lc408              :in std_logic_vector(8 DOWNTO 0);
     Lc409              :in std_logic_vector(8 DOWNTO 0);
     Lc410              :in std_logic_vector(8 DOWNTO 0);
     Lc411              :in std_logic_vector(8 DOWNTO 0);
     Lc412              :in std_logic_vector(8 DOWNTO 0);
     Lc413              :in std_logic_vector(8 DOWNTO 0);
     Lc414              :in std_logic_vector(8 DOWNTO 0);
     Lc415              :in std_logic_vector(8 DOWNTO 0);
     Lc416              :in std_logic_vector(8 DOWNTO 0);
     Lc417              :in std_logic_vector(8 DOWNTO 0);
     Lc418              :in std_logic_vector(8 DOWNTO 0);
     Lc419              :in std_logic_vector(8 DOWNTO 0);
     Lc420              :in std_logic_vector(8 DOWNTO 0);
     Lc421              :in std_logic_vector(8 DOWNTO 0);
     Lc422              :in std_logic_vector(8 DOWNTO 0);
     Lc423              :in std_logic_vector(8 DOWNTO 0);
     Lc424              :in std_logic_vector(8 DOWNTO 0);
     Lc425              :in std_logic_vector(8 DOWNTO 0);
     Lc426              :in std_logic_vector(8 DOWNTO 0);
     Lc427              :in std_logic_vector(8 DOWNTO 0);
     Lc428              :in std_logic_vector(8 DOWNTO 0);
     Lc429              :in std_logic_vector(8 DOWNTO 0);
     Lc430              :in std_logic_vector(8 DOWNTO 0);
     Lc431              :in std_logic_vector(8 DOWNTO 0);
     Lc432              :in std_logic_vector(8 DOWNTO 0);
     Lc433              :in std_logic_vector(8 DOWNTO 0);
     Lc434              :in std_logic_vector(8 DOWNTO 0);
     Lc435              :in std_logic_vector(8 DOWNTO 0);
     Lc436              :in std_logic_vector(8 DOWNTO 0);
     Lc437              :in std_logic_vector(8 DOWNTO 0);
     Lc438              :in std_logic_vector(8 DOWNTO 0);
     Lc439              :in std_logic_vector(8 DOWNTO 0);
     Lc440              :in std_logic_vector(8 DOWNTO 0);
     Lc441              :in std_logic_vector(8 DOWNTO 0);
     Lc442              :in std_logic_vector(8 DOWNTO 0);
     Lc443              :in std_logic_vector(8 DOWNTO 0);
     Lc444              :in std_logic_vector(8 DOWNTO 0);
     Lc445              :in std_logic_vector(8 DOWNTO 0);
     Lc446              :in std_logic_vector(8 DOWNTO 0);
     Lc447              :in std_logic_vector(8 DOWNTO 0);
     Lc448              :in std_logic_vector(8 DOWNTO 0);
     Lc449              :in std_logic_vector(8 DOWNTO 0);
     Lc450              :in std_logic_vector(8 DOWNTO 0);
     Lc451              :in std_logic_vector(8 DOWNTO 0);
     Lc452              :in std_logic_vector(8 DOWNTO 0);
     Lc453              :in std_logic_vector(8 DOWNTO 0);
     Lc454              :in std_logic_vector(8 DOWNTO 0);
     Lc455              :in std_logic_vector(8 DOWNTO 0);
     Lc456              :in std_logic_vector(8 DOWNTO 0);
     Lc457              :in std_logic_vector(8 DOWNTO 0);
     Lc458              :in std_logic_vector(8 DOWNTO 0);
     Lc459              :in std_logic_vector(8 DOWNTO 0);
     Lc460              :in std_logic_vector(8 DOWNTO 0);
     Lc461              :in std_logic_vector(8 DOWNTO 0);
     Lc462              :in std_logic_vector(8 DOWNTO 0);
     Lc463              :in std_logic_vector(8 DOWNTO 0);
     Lc464              :in std_logic_vector(8 DOWNTO 0);
     Lc465              :in std_logic_vector(8 DOWNTO 0);
     Lc466              :in std_logic_vector(8 DOWNTO 0);
     Lc467              :in std_logic_vector(8 DOWNTO 0);
     Lc468              :in std_logic_vector(8 DOWNTO 0);
     Lc469              :in std_logic_vector(8 DOWNTO 0);
     Lc470              :in std_logic_vector(8 DOWNTO 0);
     Lc471              :in std_logic_vector(8 DOWNTO 0);
     Lc472              :in std_logic_vector(8 DOWNTO 0);
     Lc473              :in std_logic_vector(8 DOWNTO 0);
     Lc474              :in std_logic_vector(8 DOWNTO 0);
     Lc475              :in std_logic_vector(8 DOWNTO 0);
     Lc476              :in std_logic_vector(8 DOWNTO 0);
     Lc477              :in std_logic_vector(8 DOWNTO 0);
     Lc478              :in std_logic_vector(8 DOWNTO 0);
     Lc479              :in std_logic_vector(8 DOWNTO 0);
     Lc480              :in std_logic_vector(8 DOWNTO 0);
     Lc481              :in std_logic_vector(8 DOWNTO 0);
     Lc482              :in std_logic_vector(8 DOWNTO 0);
     Lc483              :in std_logic_vector(8 DOWNTO 0);
     Lc484              :in std_logic_vector(8 DOWNTO 0);
     Lc485              :in std_logic_vector(8 DOWNTO 0);
     Lc486              :in std_logic_vector(8 DOWNTO 0);
     Lc487              :in std_logic_vector(8 DOWNTO 0);
     Lc488              :in std_logic_vector(8 DOWNTO 0);
     Lc489              :in std_logic_vector(8 DOWNTO 0);
     Lc490              :in std_logic_vector(8 DOWNTO 0);
     Lc491              :in std_logic_vector(8 DOWNTO 0);
     Lc492              :in std_logic_vector(8 DOWNTO 0);
     Lc493              :in std_logic_vector(8 DOWNTO 0);
     Lc494              :in std_logic_vector(8 DOWNTO 0);
     Lc495              :in std_logic_vector(8 DOWNTO 0);
     Lc496              :in std_logic_vector(8 DOWNTO 0);
     Lc497              :in std_logic_vector(8 DOWNTO 0);
     Lc498              :in std_logic_vector(8 DOWNTO 0);
     Lc499              :in std_logic_vector(8 DOWNTO 0);
     Lc500              :in std_logic_vector(8 DOWNTO 0);
     Lc501              :in std_logic_vector(8 DOWNTO 0);
     Lc502              :in std_logic_vector(8 DOWNTO 0);
     Lc503              :in std_logic_vector(8 DOWNTO 0);
     Lc504              :in std_logic_vector(8 DOWNTO 0);
     Lc505              :in std_logic_vector(8 DOWNTO 0);
     Lc506              :in std_logic_vector(8 DOWNTO 0);
     Lc507              :in std_logic_vector(8 DOWNTO 0);
     Lc508              :in std_logic_vector(8 DOWNTO 0);
     Lc509              :in std_logic_vector(8 DOWNTO 0);
     Lc510              :in std_logic_vector(8 DOWNTO 0);
     Lc511              :in std_logic_vector(8 DOWNTO 0);
     Lc512              :in std_logic_vector(8 DOWNTO 0);
     Lc513              :in std_logic_vector(8 DOWNTO 0);
     Lc514              :in std_logic_vector(8 DOWNTO 0);
     Lc515              :in std_logic_vector(8 DOWNTO 0);
     Lc516              :in std_logic_vector(8 DOWNTO 0);
     Lc517              :in std_logic_vector(8 DOWNTO 0);
     Lc518              :in std_logic_vector(8 DOWNTO 0);
     Lc519              :in std_logic_vector(8 DOWNTO 0);
     Lc520              :in std_logic_vector(8 DOWNTO 0);
     Lc521              :in std_logic_vector(8 DOWNTO 0);
     Lc522              :in std_logic_vector(8 DOWNTO 0);
     Lc523              :in std_logic_vector(8 DOWNTO 0);
     Lc524              :in std_logic_vector(8 DOWNTO 0);
     Lc525              :in std_logic_vector(8 DOWNTO 0);
     Lc526              :in std_logic_vector(8 DOWNTO 0);
     Lc527              :in std_logic_vector(8 DOWNTO 0);
     Lc528              :in std_logic_vector(8 DOWNTO 0);
     Lc529              :in std_logic_vector(8 DOWNTO 0);
     Lc530              :in std_logic_vector(8 DOWNTO 0);
     Lc531              :in std_logic_vector(8 DOWNTO 0);
     Lc532              :in std_logic_vector(8 DOWNTO 0);
     Lc533              :in std_logic_vector(8 DOWNTO 0);
     Lc534              :in std_logic_vector(8 DOWNTO 0);
     Lc535              :in std_logic_vector(8 DOWNTO 0);
     Lc536              :in std_logic_vector(8 DOWNTO 0);
     Lc537              :in std_logic_vector(8 DOWNTO 0);
     Lc538              :in std_logic_vector(8 DOWNTO 0);
     Lc539              :in std_logic_vector(8 DOWNTO 0);
     Lc540              :in std_logic_vector(8 DOWNTO 0);
     Lc541              :in std_logic_vector(8 DOWNTO 0);
     Lc542              :in std_logic_vector(8 DOWNTO 0);
     Lc543              :in std_logic_vector(8 DOWNTO 0);
     Lc544              :in std_logic_vector(8 DOWNTO 0);
     Lc545              :in std_logic_vector(8 DOWNTO 0);
     Lc546              :in std_logic_vector(8 DOWNTO 0);
     Lc547              :in std_logic_vector(8 DOWNTO 0);
     Lc548              :in std_logic_vector(8 DOWNTO 0);
     Lc549              :in std_logic_vector(8 DOWNTO 0);
     Lc550              :in std_logic_vector(8 DOWNTO 0);
     Lc551              :in std_logic_vector(8 DOWNTO 0);
     Lc552              :in std_logic_vector(8 DOWNTO 0);
     Lc553              :in std_logic_vector(8 DOWNTO 0);
     Lc554              :in std_logic_vector(8 DOWNTO 0);
     Lc555              :in std_logic_vector(8 DOWNTO 0);
     Lc556              :in std_logic_vector(8 DOWNTO 0);
     Lc557              :in std_logic_vector(8 DOWNTO 0);
     Lc558              :in std_logic_vector(8 DOWNTO 0);
     Lc559              :in std_logic_vector(8 DOWNTO 0);
     Lc560              :in std_logic_vector(8 DOWNTO 0);
     Lc561              :in std_logic_vector(8 DOWNTO 0);
     Lc562              :in std_logic_vector(8 DOWNTO 0);
     Lc563              :in std_logic_vector(8 DOWNTO 0);
     Lc564              :in std_logic_vector(8 DOWNTO 0);
     Lc565              :in std_logic_vector(8 DOWNTO 0);
     Lc566              :in std_logic_vector(8 DOWNTO 0);
     Lc567              :in std_logic_vector(8 DOWNTO 0);
     Lc568              :in std_logic_vector(8 DOWNTO 0);
     Lc569              :in std_logic_vector(8 DOWNTO 0);
     Lc570              :in std_logic_vector(8 DOWNTO 0);
     Lc571              :in std_logic_vector(8 DOWNTO 0);
     Lc572              :in std_logic_vector(8 DOWNTO 0);
     Lc573              :in std_logic_vector(8 DOWNTO 0);
     Lc574              :in std_logic_vector(8 DOWNTO 0);
     Lc575              :in std_logic_vector(8 DOWNTO 0);
     Lc576              :in std_logic_vector(8 DOWNTO 0);
     Lc577              :in std_logic_vector(8 DOWNTO 0);
     Lc578              :in std_logic_vector(8 DOWNTO 0);
     Lc579              :in std_logic_vector(8 DOWNTO 0);
     Lc580              :in std_logic_vector(8 DOWNTO 0);
     Lc581              :in std_logic_vector(8 DOWNTO 0);
     Lc582              :in std_logic_vector(8 DOWNTO 0);
     Lc583              :in std_logic_vector(8 DOWNTO 0);
     Lc584              :in std_logic_vector(8 DOWNTO 0);
     Lc585              :in std_logic_vector(8 DOWNTO 0);
     Lc586              :in std_logic_vector(8 DOWNTO 0);
     Lc587              :in std_logic_vector(8 DOWNTO 0);
     Lc588              :in std_logic_vector(8 DOWNTO 0);
     Lc589              :in std_logic_vector(8 DOWNTO 0);
     Lc590              :in std_logic_vector(8 DOWNTO 0);
     Lc591              :in std_logic_vector(8 DOWNTO 0);
     Lc592              :in std_logic_vector(8 DOWNTO 0);
     Lc593              :in std_logic_vector(8 DOWNTO 0);
     Lc594              :in std_logic_vector(8 DOWNTO 0);
     Lc595              :in std_logic_vector(8 DOWNTO 0);
     Lc596              :in std_logic_vector(8 DOWNTO 0);
     Lc597              :in std_logic_vector(8 DOWNTO 0);
     Lc598              :in std_logic_vector(8 DOWNTO 0);
     Lc599              :in std_logic_vector(8 DOWNTO 0);
     Lc600              :in std_logic_vector(8 DOWNTO 0);
     Lc601              :in std_logic_vector(8 DOWNTO 0);
     Lc602              :in std_logic_vector(8 DOWNTO 0);
     Lc603              :in std_logic_vector(8 DOWNTO 0);
     Lc604              :in std_logic_vector(8 DOWNTO 0);
     Lc605              :in std_logic_vector(8 DOWNTO 0);
     Lc606              :in std_logic_vector(8 DOWNTO 0);
     Lc607              :in std_logic_vector(8 DOWNTO 0);
     Lc608              :in std_logic_vector(8 DOWNTO 0);
     Lc609              :in std_logic_vector(8 DOWNTO 0);
     Lc610              :in std_logic_vector(8 DOWNTO 0);
     Lc611              :in std_logic_vector(8 DOWNTO 0);
     Lc612              :in std_logic_vector(8 DOWNTO 0);
     Lc613              :in std_logic_vector(8 DOWNTO 0);
     Lc614              :in std_logic_vector(8 DOWNTO 0);
     Lc615              :in std_logic_vector(8 DOWNTO 0);
     Lc616              :in std_logic_vector(8 DOWNTO 0);
     Lc617              :in std_logic_vector(8 DOWNTO 0);
     Lc618              :in std_logic_vector(8 DOWNTO 0);
     Lc619              :in std_logic_vector(8 DOWNTO 0);
     Lc620              :in std_logic_vector(8 DOWNTO 0);
     Lc621              :in std_logic_vector(8 DOWNTO 0);
     Lc622              :in std_logic_vector(8 DOWNTO 0);
     Lc623              :in std_logic_vector(8 DOWNTO 0);
     Lc624              :in std_logic_vector(8 DOWNTO 0);
     Lc625              :in std_logic_vector(8 DOWNTO 0);
     Lc626              :in std_logic_vector(8 DOWNTO 0);
     Lc627              :in std_logic_vector(8 DOWNTO 0);
     Lc628              :in std_logic_vector(8 DOWNTO 0);
     Lc629              :in std_logic_vector(8 DOWNTO 0);
     Lc630              :in std_logic_vector(8 DOWNTO 0);
     Lc631              :in std_logic_vector(8 DOWNTO 0);
     Lc632              :in std_logic_vector(8 DOWNTO 0);
     Lc633              :in std_logic_vector(8 DOWNTO 0);
     Lc634              :in std_logic_vector(8 DOWNTO 0);
     Lc635              :in std_logic_vector(8 DOWNTO 0);
     Lc636              :in std_logic_vector(8 DOWNTO 0);
     Lc637              :in std_logic_vector(8 DOWNTO 0);
     Lc638              :in std_logic_vector(8 DOWNTO 0);
     Lc639              :in std_logic_vector(8 DOWNTO 0);
     Lc640              :in std_logic_vector(8 DOWNTO 0);
     Lc641              :in std_logic_vector(8 DOWNTO 0);
     Lc642              :in std_logic_vector(8 DOWNTO 0);
     Lc643              :in std_logic_vector(8 DOWNTO 0);
     Lc644              :in std_logic_vector(8 DOWNTO 0);
     Lc645              :in std_logic_vector(8 DOWNTO 0);
     Lc646              :in std_logic_vector(8 DOWNTO 0);
     Lc647              :in std_logic_vector(8 DOWNTO 0);
     Lc648              :in std_logic_vector(8 DOWNTO 0);
     Lc649              :in std_logic_vector(8 DOWNTO 0);
     Lc650              :in std_logic_vector(8 DOWNTO 0);
     Lc651              :in std_logic_vector(8 DOWNTO 0);
     Lc652              :in std_logic_vector(8 DOWNTO 0);
     Lc653              :in std_logic_vector(8 DOWNTO 0);
     Lc654              :in std_logic_vector(8 DOWNTO 0);
     Lc655              :in std_logic_vector(8 DOWNTO 0);
     Lc656              :in std_logic_vector(8 DOWNTO 0);
     Lc657              :in std_logic_vector(8 DOWNTO 0);
     Lc658              :in std_logic_vector(8 DOWNTO 0);
     Lc659              :in std_logic_vector(8 DOWNTO 0);
     Lc660              :in std_logic_vector(8 DOWNTO 0);
     Lc661              :in std_logic_vector(8 DOWNTO 0);
     Lc662              :in std_logic_vector(8 DOWNTO 0);
     Lc663              :in std_logic_vector(8 DOWNTO 0);
     Lc664              :in std_logic_vector(8 DOWNTO 0);
     Lc665              :in std_logic_vector(8 DOWNTO 0);
     Lc666              :in std_logic_vector(8 DOWNTO 0);
     Lc667              :in std_logic_vector(8 DOWNTO 0);
     Lc668              :in std_logic_vector(8 DOWNTO 0);
     Lc669              :in std_logic_vector(8 DOWNTO 0);
     Lc670              :in std_logic_vector(8 DOWNTO 0);
     Lc671              :in std_logic_vector(8 DOWNTO 0);
     Lc672              :in std_logic_vector(8 DOWNTO 0);
     Lc673              :in std_logic_vector(8 DOWNTO 0);
     Lc674              :in std_logic_vector(8 DOWNTO 0);
     Lc675              :in std_logic_vector(8 DOWNTO 0);
     Lc676              :in std_logic_vector(8 DOWNTO 0);
     Lc677              :in std_logic_vector(8 DOWNTO 0);
     Lc678              :in std_logic_vector(8 DOWNTO 0);
     Lc679              :in std_logic_vector(8 DOWNTO 0);
     Lc680              :in std_logic_vector(8 DOWNTO 0);
     Lc681              :in std_logic_vector(8 DOWNTO 0);
     Lc682              :in std_logic_vector(8 DOWNTO 0);
     Lc683              :in std_logic_vector(8 DOWNTO 0);
     Lc684              :in std_logic_vector(8 DOWNTO 0);
     Lc685              :in std_logic_vector(8 DOWNTO 0);
     Lc686              :in std_logic_vector(8 DOWNTO 0);
     Lc687              :in std_logic_vector(8 DOWNTO 0);
     Lc688              :in std_logic_vector(8 DOWNTO 0);
     Lc689              :in std_logic_vector(8 DOWNTO 0);
     Lc690              :in std_logic_vector(8 DOWNTO 0);
     Lc691              :in std_logic_vector(8 DOWNTO 0);
     Lc692              :in std_logic_vector(8 DOWNTO 0);
     Lc693              :in std_logic_vector(8 DOWNTO 0);
     Lc694              :in std_logic_vector(8 DOWNTO 0);
     Lc695              :in std_logic_vector(8 DOWNTO 0);
     Lc696              :in std_logic_vector(8 DOWNTO 0);
     Lc697              :in std_logic_vector(8 DOWNTO 0);
     Lc698              :in std_logic_vector(8 DOWNTO 0);
     Lc699              :in std_logic_vector(8 DOWNTO 0);
     Lc700              :in std_logic_vector(8 DOWNTO 0);
     Lc701              :in std_logic_vector(8 DOWNTO 0);
     Lc702              :in std_logic_vector(8 DOWNTO 0);
     Lc703              :in std_logic_vector(8 DOWNTO 0);
     Lc704              :in std_logic_vector(8 DOWNTO 0);
     Lc705              :in std_logic_vector(8 DOWNTO 0);
     Lc706              :in std_logic_vector(8 DOWNTO 0);
     Lc707              :in std_logic_vector(8 DOWNTO 0);
     Lc708              :in std_logic_vector(8 DOWNTO 0);
     Lc709              :in std_logic_vector(8 DOWNTO 0);
     Lc710              :in std_logic_vector(8 DOWNTO 0);
     Lc711              :in std_logic_vector(8 DOWNTO 0);
     Lc712              :in std_logic_vector(8 DOWNTO 0);
     Lc713              :in std_logic_vector(8 DOWNTO 0);
     Lc714              :in std_logic_vector(8 DOWNTO 0);
     Lc715              :in std_logic_vector(8 DOWNTO 0);
     Lc716              :in std_logic_vector(8 DOWNTO 0);
     Lc717              :in std_logic_vector(8 DOWNTO 0);
     Lc718              :in std_logic_vector(8 DOWNTO 0);
     Lc719              :in std_logic_vector(8 DOWNTO 0);
     Lc720              :in std_logic_vector(8 DOWNTO 0);
     Lc721              :in std_logic_vector(8 DOWNTO 0);
     Lc722              :in std_logic_vector(8 DOWNTO 0);
     Lc723              :in std_logic_vector(8 DOWNTO 0);
     Lc724              :in std_logic_vector(8 DOWNTO 0);
     Lc725              :in std_logic_vector(8 DOWNTO 0);
     Lc726              :in std_logic_vector(8 DOWNTO 0);
     Lc727              :in std_logic_vector(8 DOWNTO 0);
     Lc728              :in std_logic_vector(8 DOWNTO 0);
     Lc729              :in std_logic_vector(8 DOWNTO 0);
     Lc730              :in std_logic_vector(8 DOWNTO 0);
     Lc731              :in std_logic_vector(8 DOWNTO 0);
     Lc732              :in std_logic_vector(8 DOWNTO 0);
     Lc733              :in std_logic_vector(8 DOWNTO 0);
     Lc734              :in std_logic_vector(8 DOWNTO 0);
     Lc735              :in std_logic_vector(8 DOWNTO 0);
     Lc736              :in std_logic_vector(8 DOWNTO 0);
     Lc737              :in std_logic_vector(8 DOWNTO 0);
     Lc738              :in std_logic_vector(8 DOWNTO 0);
     Lc739              :in std_logic_vector(8 DOWNTO 0);
     Lc740              :in std_logic_vector(8 DOWNTO 0);
     Lc741              :in std_logic_vector(8 DOWNTO 0);
     Lc742              :in std_logic_vector(8 DOWNTO 0);
     Lc743              :in std_logic_vector(8 DOWNTO 0);
     Lc744              :in std_logic_vector(8 DOWNTO 0);
     Lc745              :in std_logic_vector(8 DOWNTO 0);
     Lc746              :in std_logic_vector(8 DOWNTO 0);
     Lc747              :in std_logic_vector(8 DOWNTO 0);
     Lc748              :in std_logic_vector(8 DOWNTO 0);
     Lc749              :in std_logic_vector(8 DOWNTO 0);
     Lc750              :in std_logic_vector(8 DOWNTO 0);
     Lc751              :in std_logic_vector(8 DOWNTO 0);
     Lc752              :in std_logic_vector(8 DOWNTO 0);
     Lc753              :in std_logic_vector(8 DOWNTO 0);
     Lc754              :in std_logic_vector(8 DOWNTO 0);
     Lc755              :in std_logic_vector(8 DOWNTO 0);
     Lc756              :in std_logic_vector(8 DOWNTO 0);
     Lc757              :in std_logic_vector(8 DOWNTO 0);
     Lc758              :in std_logic_vector(8 DOWNTO 0);
     Lc759              :in std_logic_vector(8 DOWNTO 0);
     Lc760              :in std_logic_vector(8 DOWNTO 0);
     Lc761              :in std_logic_vector(8 DOWNTO 0);
     Lc762              :in std_logic_vector(8 DOWNTO 0);
     Lc763              :in std_logic_vector(8 DOWNTO 0);
     Lc764              :in std_logic_vector(8 DOWNTO 0);
     Lc765              :in std_logic_vector(8 DOWNTO 0);
     Lc766              :in std_logic_vector(8 DOWNTO 0);
     Lc767              :in std_logic_vector(8 DOWNTO 0);
     Lc768              :in std_logic_vector(8 DOWNTO 0);
     Lc769              :in std_logic_vector(8 DOWNTO 0);
     Lc770              :in std_logic_vector(8 DOWNTO 0);
     Lc771              :in std_logic_vector(8 DOWNTO 0);
     Lc772              :in std_logic_vector(8 DOWNTO 0);
     Lc773              :in std_logic_vector(8 DOWNTO 0);
     Lc774              :in std_logic_vector(8 DOWNTO 0);
     Lc775              :in std_logic_vector(8 DOWNTO 0);
     Lc776              :in std_logic_vector(8 DOWNTO 0);
     Lc777              :in std_logic_vector(8 DOWNTO 0);
     Lc778              :in std_logic_vector(8 DOWNTO 0);
     Lc779              :in std_logic_vector(8 DOWNTO 0);
     Lc780              :in std_logic_vector(8 DOWNTO 0);
     Lc781              :in std_logic_vector(8 DOWNTO 0);
     Lc782              :in std_logic_vector(8 DOWNTO 0);
     Lc783              :in std_logic_vector(8 DOWNTO 0);
     Lc784              :in std_logic_vector(8 DOWNTO 0);
     Lc785              :in std_logic_vector(8 DOWNTO 0);
     Lc786              :in std_logic_vector(8 DOWNTO 0);
     Lc787              :in std_logic_vector(8 DOWNTO 0);
     Lc788              :in std_logic_vector(8 DOWNTO 0);
     Lc789              :in std_logic_vector(8 DOWNTO 0);
     Lc790              :in std_logic_vector(8 DOWNTO 0);
     Lc791              :in std_logic_vector(8 DOWNTO 0);
     Lc792              :in std_logic_vector(8 DOWNTO 0);
     Lc793              :in std_logic_vector(8 DOWNTO 0);
     Lc794              :in std_logic_vector(8 DOWNTO 0);
     Lc795              :in std_logic_vector(8 DOWNTO 0);
     Lc796              :in std_logic_vector(8 DOWNTO 0);
     Lc797              :in std_logic_vector(8 DOWNTO 0);
     Lc798              :in std_logic_vector(8 DOWNTO 0);
     Lc799              :in std_logic_vector(8 DOWNTO 0);
     Lc800              :in std_logic_vector(8 DOWNTO 0);
     Lc801              :in std_logic_vector(8 DOWNTO 0);
     Lc802              :in std_logic_vector(8 DOWNTO 0);
     Lc803              :in std_logic_vector(8 DOWNTO 0);
     Lc804              :in std_logic_vector(8 DOWNTO 0);
     Lc805              :in std_logic_vector(8 DOWNTO 0);
     Lc806              :in std_logic_vector(8 DOWNTO 0);
     Lc807              :in std_logic_vector(8 DOWNTO 0);
     Lc808              :in std_logic_vector(8 DOWNTO 0);
     Lc809              :in std_logic_vector(8 DOWNTO 0);
     Lc810              :in std_logic_vector(8 DOWNTO 0);
     Lc811              :in std_logic_vector(8 DOWNTO 0);
     Lc812              :in std_logic_vector(8 DOWNTO 0);
     Lc813              :in std_logic_vector(8 DOWNTO 0);
     Lc814              :in std_logic_vector(8 DOWNTO 0);
     Lc815              :in std_logic_vector(8 DOWNTO 0);
     Lc816              :in std_logic_vector(8 DOWNTO 0);
     Lc817              :in std_logic_vector(8 DOWNTO 0);
     Lc818              :in std_logic_vector(8 DOWNTO 0);
     Lc819              :in std_logic_vector(8 DOWNTO 0);
     Lc820              :in std_logic_vector(8 DOWNTO 0);
     Lc821              :in std_logic_vector(8 DOWNTO 0);
     Lc822              :in std_logic_vector(8 DOWNTO 0);
     Lc823              :in std_logic_vector(8 DOWNTO 0);
     Lc824              :in std_logic_vector(8 DOWNTO 0);
     Lc825              :in std_logic_vector(8 DOWNTO 0);
     Lc826              :in std_logic_vector(8 DOWNTO 0);
     Lc827              :in std_logic_vector(8 DOWNTO 0);
     Lc828              :in std_logic_vector(8 DOWNTO 0);
     Lc829              :in std_logic_vector(8 DOWNTO 0);
     Lc830              :in std_logic_vector(8 DOWNTO 0);
     Lc831              :in std_logic_vector(8 DOWNTO 0);
     Lc832              :in std_logic_vector(8 DOWNTO 0);
     Lc833              :in std_logic_vector(8 DOWNTO 0);
     Lc834              :in std_logic_vector(8 DOWNTO 0);
     Lc835              :in std_logic_vector(8 DOWNTO 0);
     Lc836              :in std_logic_vector(8 DOWNTO 0);
     Lc837              :in std_logic_vector(8 DOWNTO 0);
     Lc838              :in std_logic_vector(8 DOWNTO 0);
     Lc839              :in std_logic_vector(8 DOWNTO 0);
     Lc840              :in std_logic_vector(8 DOWNTO 0);
     Lc841              :in std_logic_vector(8 DOWNTO 0);
     Lc842              :in std_logic_vector(8 DOWNTO 0);
     Lc843              :in std_logic_vector(8 DOWNTO 0);
     Lc844              :in std_logic_vector(8 DOWNTO 0);
     Lc845              :in std_logic_vector(8 DOWNTO 0);
     Lc846              :in std_logic_vector(8 DOWNTO 0);
     Lc847              :in std_logic_vector(8 DOWNTO 0);
     Lc848              :in std_logic_vector(8 DOWNTO 0);
     Lc849              :in std_logic_vector(8 DOWNTO 0);
     Lc850              :in std_logic_vector(8 DOWNTO 0);
     Lc851              :in std_logic_vector(8 DOWNTO 0);
     Lc852              :in std_logic_vector(8 DOWNTO 0);
     Lc853              :in std_logic_vector(8 DOWNTO 0);
     Lc854              :in std_logic_vector(8 DOWNTO 0);
     Lc855              :in std_logic_vector(8 DOWNTO 0);
     Lc856              :in std_logic_vector(8 DOWNTO 0);
     Lc857              :in std_logic_vector(8 DOWNTO 0);
     Lc858              :in std_logic_vector(8 DOWNTO 0);
     Lc859              :in std_logic_vector(8 DOWNTO 0);
     Lc860              :in std_logic_vector(8 DOWNTO 0);
     Lc861              :in std_logic_vector(8 DOWNTO 0);
     Lc862              :in std_logic_vector(8 DOWNTO 0);
     Lc863              :in std_logic_vector(8 DOWNTO 0);
     Lc864              :in std_logic_vector(8 DOWNTO 0);
     Lc865              :in std_logic_vector(8 DOWNTO 0);
     Lc866              :in std_logic_vector(8 DOWNTO 0);
     Lc867              :in std_logic_vector(8 DOWNTO 0);
     Lc868              :in std_logic_vector(8 DOWNTO 0);
     Lc869              :in std_logic_vector(8 DOWNTO 0);
     Lc870              :in std_logic_vector(8 DOWNTO 0);
     Lc871              :in std_logic_vector(8 DOWNTO 0);
     Lc872              :in std_logic_vector(8 DOWNTO 0);
     Lc873              :in std_logic_vector(8 DOWNTO 0);
     Lc874              :in std_logic_vector(8 DOWNTO 0);
     Lc875              :in std_logic_vector(8 DOWNTO 0);
     Lc876              :in std_logic_vector(8 DOWNTO 0);
     Lc877              :in std_logic_vector(8 DOWNTO 0);
     Lc878              :in std_logic_vector(8 DOWNTO 0);
     Lc879              :in std_logic_vector(8 DOWNTO 0);
     Lc880              :in std_logic_vector(8 DOWNTO 0);
     Lc881              :in std_logic_vector(8 DOWNTO 0);
     Lc882              :in std_logic_vector(8 DOWNTO 0);
     Lc883              :in std_logic_vector(8 DOWNTO 0);
     Lc884              :in std_logic_vector(8 DOWNTO 0);
     Lc885              :in std_logic_vector(8 DOWNTO 0);
     Lc886              :in std_logic_vector(8 DOWNTO 0);
     Lc887              :in std_logic_vector(8 DOWNTO 0);
     Lc888              :in std_logic_vector(8 DOWNTO 0);
     Lc889              :in std_logic_vector(8 DOWNTO 0);
     Lc890              :in std_logic_vector(8 DOWNTO 0);
     Lc891              :in std_logic_vector(8 DOWNTO 0);
     Lc892              :in std_logic_vector(8 DOWNTO 0);
     Lc893              :in std_logic_vector(8 DOWNTO 0);
     Lc894              :in std_logic_vector(8 DOWNTO 0);
     Lc895              :in std_logic_vector(8 DOWNTO 0);
     Lc896              :in std_logic_vector(8 DOWNTO 0);
     Lc897              :in std_logic_vector(8 DOWNTO 0);
     Lc898              :in std_logic_vector(8 DOWNTO 0);
     Lc899              :in std_logic_vector(8 DOWNTO 0);
     Lc900              :in std_logic_vector(8 DOWNTO 0);
     Lc901              :in std_logic_vector(8 DOWNTO 0);
     Lc902              :in std_logic_vector(8 DOWNTO 0);
     Lc903              :in std_logic_vector(8 DOWNTO 0);
     Lc904              :in std_logic_vector(8 DOWNTO 0);
     Lc905              :in std_logic_vector(8 DOWNTO 0);
     Lc906              :in std_logic_vector(8 DOWNTO 0);
     Lc907              :in std_logic_vector(8 DOWNTO 0);
     Lc908              :in std_logic_vector(8 DOWNTO 0);
     Lc909              :in std_logic_vector(8 DOWNTO 0);
     Lc910              :in std_logic_vector(8 DOWNTO 0);
     Lc911              :in std_logic_vector(8 DOWNTO 0);
     Lc912              :in std_logic_vector(8 DOWNTO 0);
     Lc913              :in std_logic_vector(8 DOWNTO 0);
     Lc914              :in std_logic_vector(8 DOWNTO 0);
     Lc915              :in std_logic_vector(8 DOWNTO 0);
     Lc916              :in std_logic_vector(8 DOWNTO 0);
     Lc917              :in std_logic_vector(8 DOWNTO 0);
     Lc918              :in std_logic_vector(8 DOWNTO 0);
     Lc919              :in std_logic_vector(8 DOWNTO 0);
     Lc920              :in std_logic_vector(8 DOWNTO 0);
     Lc921              :in std_logic_vector(8 DOWNTO 0);
     Lc922              :in std_logic_vector(8 DOWNTO 0);
     Lc923              :in std_logic_vector(8 DOWNTO 0);
     Lc924              :in std_logic_vector(8 DOWNTO 0);
     Lc925              :in std_logic_vector(8 DOWNTO 0);
     Lc926              :in std_logic_vector(8 DOWNTO 0);
     Lc927              :in std_logic_vector(8 DOWNTO 0);
     Lc928              :in std_logic_vector(8 DOWNTO 0);
     Lc929              :in std_logic_vector(8 DOWNTO 0);
     Lc930              :in std_logic_vector(8 DOWNTO 0);
     Lc931              :in std_logic_vector(8 DOWNTO 0);
     Lc932              :in std_logic_vector(8 DOWNTO 0);
     Lc933              :in std_logic_vector(8 DOWNTO 0);
     Lc934              :in std_logic_vector(8 DOWNTO 0);
     Lc935              :in std_logic_vector(8 DOWNTO 0);
     Lc936              :in std_logic_vector(8 DOWNTO 0);
     Lc937              :in std_logic_vector(8 DOWNTO 0);
     Lc938              :in std_logic_vector(8 DOWNTO 0);
     Lc939              :in std_logic_vector(8 DOWNTO 0);
     Lc940              :in std_logic_vector(8 DOWNTO 0);
     Lc941              :in std_logic_vector(8 DOWNTO 0);
     Lc942              :in std_logic_vector(8 DOWNTO 0);
     Lc943              :in std_logic_vector(8 DOWNTO 0);
     Lc944              :in std_logic_vector(8 DOWNTO 0);
     Lc945              :in std_logic_vector(8 DOWNTO 0);
     Lc946              :in std_logic_vector(8 DOWNTO 0);
     Lc947              :in std_logic_vector(8 DOWNTO 0);
     Lc948              :in std_logic_vector(8 DOWNTO 0);
     Lc949              :in std_logic_vector(8 DOWNTO 0);
     Lc950              :in std_logic_vector(8 DOWNTO 0);
     Lc951              :in std_logic_vector(8 DOWNTO 0);
     Lc952              :in std_logic_vector(8 DOWNTO 0);
     Lc953              :in std_logic_vector(8 DOWNTO 0);
     Lc954              :in std_logic_vector(8 DOWNTO 0);
     Lc955              :in std_logic_vector(8 DOWNTO 0);
     Lc956              :in std_logic_vector(8 DOWNTO 0);
     Lc957              :in std_logic_vector(8 DOWNTO 0);
     Lc958              :in std_logic_vector(8 DOWNTO 0);
     Lc959              :in std_logic_vector(8 DOWNTO 0);
     Lc960              :in std_logic_vector(8 DOWNTO 0);
     Lc961              :in std_logic_vector(8 DOWNTO 0);
     Lc962              :in std_logic_vector(8 DOWNTO 0);
     Lc963              :in std_logic_vector(8 DOWNTO 0);
     Lc964              :in std_logic_vector(8 DOWNTO 0);
     Lc965              :in std_logic_vector(8 DOWNTO 0);
     Lc966              :in std_logic_vector(8 DOWNTO 0);
     Lc967              :in std_logic_vector(8 DOWNTO 0);
     Lc968              :in std_logic_vector(8 DOWNTO 0);
     Lc969              :in std_logic_vector(8 DOWNTO 0);
     Lc970              :in std_logic_vector(8 DOWNTO 0);
     Lc971              :in std_logic_vector(8 DOWNTO 0);
     Lc972              :in std_logic_vector(8 DOWNTO 0);
     Lc973              :in std_logic_vector(8 DOWNTO 0);
     Lc974              :in std_logic_vector(8 DOWNTO 0);
     Lc975              :in std_logic_vector(8 DOWNTO 0);
     Lc976              :in std_logic_vector(8 DOWNTO 0);
     Lc977              :in std_logic_vector(8 DOWNTO 0);
     Lc978              :in std_logic_vector(8 DOWNTO 0);
     Lc979              :in std_logic_vector(8 DOWNTO 0);
     Lc980              :in std_logic_vector(8 DOWNTO 0);
     Lc981              :in std_logic_vector(8 DOWNTO 0);
     Lc982              :in std_logic_vector(8 DOWNTO 0);
     Lc983              :in std_logic_vector(8 DOWNTO 0);
     Lc984              :in std_logic_vector(8 DOWNTO 0);
     Lc985              :in std_logic_vector(8 DOWNTO 0);
     Lc986              :in std_logic_vector(8 DOWNTO 0);
     Lc987              :in std_logic_vector(8 DOWNTO 0);
     Lc988              :in std_logic_vector(8 DOWNTO 0);
     Lc989              :in std_logic_vector(8 DOWNTO 0);
     Lc990              :in std_logic_vector(8 DOWNTO 0);
     Lc991              :in std_logic_vector(8 DOWNTO 0);
     Lc992              :in std_logic_vector(8 DOWNTO 0);
     Lc993              :in std_logic_vector(8 DOWNTO 0);
     Lc994              :in std_logic_vector(8 DOWNTO 0);
     Lc995              :in std_logic_vector(8 DOWNTO 0);
     Lc996              :in std_logic_vector(8 DOWNTO 0);
     Lc997              :in std_logic_vector(8 DOWNTO 0);
     Lc998              :in std_logic_vector(8 DOWNTO 0);
     Lc999              :in std_logic_vector(8 DOWNTO 0);
     Lc1000              :in std_logic_vector(8 DOWNTO 0);
     Lc1001              :in std_logic_vector(8 DOWNTO 0);
     Lc1002              :in std_logic_vector(8 DOWNTO 0);
     Lc1003              :in std_logic_vector(8 DOWNTO 0);
     Lc1004              :in std_logic_vector(8 DOWNTO 0);
     Lc1005              :in std_logic_vector(8 DOWNTO 0);
     Lc1006              :in std_logic_vector(8 DOWNTO 0);
     Lc1007              :in std_logic_vector(8 DOWNTO 0);
     Lc1008              :in std_logic_vector(8 DOWNTO 0);
     Lc1009              :in std_logic_vector(8 DOWNTO 0);
     Lc1010              :in std_logic_vector(8 DOWNTO 0);
     Lc1011              :in std_logic_vector(8 DOWNTO 0);
     Lc1012              :in std_logic_vector(8 DOWNTO 0);
     Lc1013              :in std_logic_vector(8 DOWNTO 0);
     Lc1014              :in std_logic_vector(8 DOWNTO 0);
     Lc1015              :in std_logic_vector(8 DOWNTO 0);
     Lc1016              :in std_logic_vector(8 DOWNTO 0);
     Lc1017              :in std_logic_vector(8 DOWNTO 0);
     Lc1018              :in std_logic_vector(8 DOWNTO 0);
     Lc1019              :in std_logic_vector(8 DOWNTO 0);
     Lc1020              :in std_logic_vector(8 DOWNTO 0);
     Lc1021              :in std_logic_vector(8 DOWNTO 0);
     Lc1022              :in std_logic_vector(8 DOWNTO 0);
     Lc1023              :in std_logic_vector(8 DOWNTO 0);
     Lc1024              :in std_logic_vector(8 DOWNTO 0);
     Lc1025              :in std_logic_vector(8 DOWNTO 0);
     Lc1026              :in std_logic_vector(8 DOWNTO 0);
     Lc1027              :in std_logic_vector(8 DOWNTO 0);
     Lc1028              :in std_logic_vector(8 DOWNTO 0);
     Lc1029              :in std_logic_vector(8 DOWNTO 0);
     Lc1030              :in std_logic_vector(8 DOWNTO 0);
     Lc1031              :in std_logic_vector(8 DOWNTO 0);
     Lc1032              :in std_logic_vector(8 DOWNTO 0);
     Lc1033              :in std_logic_vector(8 DOWNTO 0);
     Lc1034              :in std_logic_vector(8 DOWNTO 0);
     Lc1035              :in std_logic_vector(8 DOWNTO 0);
     Lc1036              :in std_logic_vector(8 DOWNTO 0);
     Lc1037              :in std_logic_vector(8 DOWNTO 0);
     Lc1038              :in std_logic_vector(8 DOWNTO 0);
     Lc1039              :in std_logic_vector(8 DOWNTO 0);
     Lc1040              :in std_logic_vector(8 DOWNTO 0);
     Lc1041              :in std_logic_vector(8 DOWNTO 0);
     Lc1042              :in std_logic_vector(8 DOWNTO 0);
     Lc1043              :in std_logic_vector(8 DOWNTO 0);
     Lc1044              :in std_logic_vector(8 DOWNTO 0);
     Lc1045              :in std_logic_vector(8 DOWNTO 0);
     Lc1046              :in std_logic_vector(8 DOWNTO 0);
     Lc1047              :in std_logic_vector(8 DOWNTO 0);
     Lc1048              :in std_logic_vector(8 DOWNTO 0);
     Lc1049              :in std_logic_vector(8 DOWNTO 0);
     Lc1050              :in std_logic_vector(8 DOWNTO 0);
     Lc1051              :in std_logic_vector(8 DOWNTO 0);
     Lc1052              :in std_logic_vector(8 DOWNTO 0);
     Lc1053              :in std_logic_vector(8 DOWNTO 0);
     Lc1054              :in std_logic_vector(8 DOWNTO 0);
     Lc1055              :in std_logic_vector(8 DOWNTO 0);
     Lc1056              :in std_logic_vector(8 DOWNTO 0);
     Lc1057              :in std_logic_vector(8 DOWNTO 0);
     Lc1058              :in std_logic_vector(8 DOWNTO 0);
     Lc1059              :in std_logic_vector(8 DOWNTO 0);
     Lc1060              :in std_logic_vector(8 DOWNTO 0);
     Lc1061              :in std_logic_vector(8 DOWNTO 0);
     Lc1062              :in std_logic_vector(8 DOWNTO 0);
     Lc1063              :in std_logic_vector(8 DOWNTO 0);
     Lc1064              :in std_logic_vector(8 DOWNTO 0);
     Lc1065              :in std_logic_vector(8 DOWNTO 0);
     Lc1066              :in std_logic_vector(8 DOWNTO 0);
     Lc1067              :in std_logic_vector(8 DOWNTO 0);
     Lc1068              :in std_logic_vector(8 DOWNTO 0);
     Lc1069              :in std_logic_vector(8 DOWNTO 0);
     Lc1070              :in std_logic_vector(8 DOWNTO 0);
     Lc1071              :in std_logic_vector(8 DOWNTO 0);
     Lc1072              :in std_logic_vector(8 DOWNTO 0);
     Lc1073              :in std_logic_vector(8 DOWNTO 0);
     Lc1074              :in std_logic_vector(8 DOWNTO 0);
     Lc1075              :in std_logic_vector(8 DOWNTO 0);
     Lc1076              :in std_logic_vector(8 DOWNTO 0);
     Lc1077              :in std_logic_vector(8 DOWNTO 0);
     Lc1078              :in std_logic_vector(8 DOWNTO 0);
     Lc1079              :in std_logic_vector(8 DOWNTO 0);
     Lc1080              :in std_logic_vector(8 DOWNTO 0);
     Lc1081              :in std_logic_vector(8 DOWNTO 0);
     Lc1082              :in std_logic_vector(8 DOWNTO 0);
     Lc1083              :in std_logic_vector(8 DOWNTO 0);
     Lc1084              :in std_logic_vector(8 DOWNTO 0);
     Lc1085              :in std_logic_vector(8 DOWNTO 0);
     Lc1086              :in std_logic_vector(8 DOWNTO 0);
     Lc1087              :in std_logic_vector(8 DOWNTO 0);
     Lc1088              :in std_logic_vector(8 DOWNTO 0);
     Lc1089              :in std_logic_vector(8 DOWNTO 0);
     Lc1090              :in std_logic_vector(8 DOWNTO 0);
     Lc1091              :in std_logic_vector(8 DOWNTO 0);
     Lc1092              :in std_logic_vector(8 DOWNTO 0);
     Lc1093              :in std_logic_vector(8 DOWNTO 0);
     Lc1094              :in std_logic_vector(8 DOWNTO 0);
     Lc1095              :in std_logic_vector(8 DOWNTO 0);
     Lc1096              :in std_logic_vector(8 DOWNTO 0);
     Lc1097              :in std_logic_vector(8 DOWNTO 0);
     Lc1098              :in std_logic_vector(8 DOWNTO 0);
     Lc1099              :in std_logic_vector(8 DOWNTO 0);
     Lc1100              :in std_logic_vector(8 DOWNTO 0);
     Lc1101              :in std_logic_vector(8 DOWNTO 0);
     Lc1102              :in std_logic_vector(8 DOWNTO 0);
     Lc1103              :in std_logic_vector(8 DOWNTO 0);
     Lc1104              :in std_logic_vector(8 DOWNTO 0);
     Lc1105              :in std_logic_vector(8 DOWNTO 0);
     Lc1106              :in std_logic_vector(8 DOWNTO 0);
     Lc1107              :in std_logic_vector(8 DOWNTO 0);
     Lc1108              :in std_logic_vector(8 DOWNTO 0);
     Lc1109              :in std_logic_vector(8 DOWNTO 0);
     Lc1110              :in std_logic_vector(8 DOWNTO 0);
     Lc1111              :in std_logic_vector(8 DOWNTO 0);
     Lc1112              :in std_logic_vector(8 DOWNTO 0);
     Lc1113              :in std_logic_vector(8 DOWNTO 0);
     Lc1114              :in std_logic_vector(8 DOWNTO 0);
     Lc1115              :in std_logic_vector(8 DOWNTO 0);
     Lc1116              :in std_logic_vector(8 DOWNTO 0);
     Lc1117              :in std_logic_vector(8 DOWNTO 0);
     Lc1118              :in std_logic_vector(8 DOWNTO 0);
     Lc1119              :in std_logic_vector(8 DOWNTO 0);
     Lc1120              :in std_logic_vector(8 DOWNTO 0);
     Lc1121              :in std_logic_vector(8 DOWNTO 0);
     Lc1122              :in std_logic_vector(8 DOWNTO 0);
     Lc1123              :in std_logic_vector(8 DOWNTO 0);
     Lc1124              :in std_logic_vector(8 DOWNTO 0);
     Lc1125              :in std_logic_vector(8 DOWNTO 0);
     Lc1126              :in std_logic_vector(8 DOWNTO 0);
     Lc1127              :in std_logic_vector(8 DOWNTO 0);
     Lc1128              :in std_logic_vector(8 DOWNTO 0);
     Lc1129              :in std_logic_vector(8 DOWNTO 0);
     Lc1130              :in std_logic_vector(8 DOWNTO 0);
     Lc1131              :in std_logic_vector(8 DOWNTO 0);
     Lc1132              :in std_logic_vector(8 DOWNTO 0);
     Lc1133              :in std_logic_vector(8 DOWNTO 0);
     Lc1134              :in std_logic_vector(8 DOWNTO 0);
     Lc1135              :in std_logic_vector(8 DOWNTO 0);
     Lc1136              :in std_logic_vector(8 DOWNTO 0);
     Lc1137              :in std_logic_vector(8 DOWNTO 0);
     Lc1138              :in std_logic_vector(8 DOWNTO 0);
     Lc1139              :in std_logic_vector(8 DOWNTO 0);
     Lc1140              :in std_logic_vector(8 DOWNTO 0);
     Lc1141              :in std_logic_vector(8 DOWNTO 0);
     Lc1142              :in std_logic_vector(8 DOWNTO 0);
     Lc1143              :in std_logic_vector(8 DOWNTO 0);
     Lc1144              :in std_logic_vector(8 DOWNTO 0);
     Lc1145              :in std_logic_vector(8 DOWNTO 0);
     Lc1146              :in std_logic_vector(8 DOWNTO 0);
     Lc1147              :in std_logic_vector(8 DOWNTO 0);
     Lc1148              :in std_logic_vector(8 DOWNTO 0);
     Lc1149              :in std_logic_vector(8 DOWNTO 0);
     Lc1150              :in std_logic_vector(8 DOWNTO 0);
     Lc1151              :in std_logic_vector(8 DOWNTO 0);
     Lc1152              :in std_logic_vector(8 DOWNTO 0);
     Lc1153              :in std_logic_vector(8 DOWNTO 0);
     Lc1154              :in std_logic_vector(8 DOWNTO 0);
     Lc1155              :in std_logic_vector(8 DOWNTO 0);
     Lc1156              :in std_logic_vector(8 DOWNTO 0);
     Lc1157              :in std_logic_vector(8 DOWNTO 0);
     Lc1158              :in std_logic_vector(8 DOWNTO 0);
     Lc1159              :in std_logic_vector(8 DOWNTO 0);
     Lc1160              :in std_logic_vector(8 DOWNTO 0);
     Lc1161              :in std_logic_vector(8 DOWNTO 0);
     Lc1162              :in std_logic_vector(8 DOWNTO 0);
     Lc1163              :in std_logic_vector(8 DOWNTO 0);
     Lc1164              :in std_logic_vector(8 DOWNTO 0);
     Lc1165              :in std_logic_vector(8 DOWNTO 0);
     Lc1166              :in std_logic_vector(8 DOWNTO 0);
     Lc1167              :in std_logic_vector(8 DOWNTO 0);
     Lc1168              :in std_logic_vector(8 DOWNTO 0);
     Lc1169              :in std_logic_vector(8 DOWNTO 0);
     Lc1170              :in std_logic_vector(8 DOWNTO 0);
     Lc1171              :in std_logic_vector(8 DOWNTO 0);
     Lc1172              :in std_logic_vector(8 DOWNTO 0);
     Lc1173              :in std_logic_vector(8 DOWNTO 0);
     Lc1174              :in std_logic_vector(8 DOWNTO 0);
     Lc1175              :in std_logic_vector(8 DOWNTO 0);
     Lc1176              :in std_logic_vector(8 DOWNTO 0);
     Lc1177              :in std_logic_vector(8 DOWNTO 0);
     Lc1178              :in std_logic_vector(8 DOWNTO 0);
     Lc1179              :in std_logic_vector(8 DOWNTO 0);
     Lc1180              :in std_logic_vector(8 DOWNTO 0);
     Lc1181              :in std_logic_vector(8 DOWNTO 0);
     Lc1182              :in std_logic_vector(8 DOWNTO 0);
     Lc1183              :in std_logic_vector(8 DOWNTO 0);
     Lc1184              :in std_logic_vector(8 DOWNTO 0);
     Lc1185              :in std_logic_vector(8 DOWNTO 0);
     Lc1186              :in std_logic_vector(8 DOWNTO 0);
     Lc1187              :in std_logic_vector(8 DOWNTO 0);
     Lc1188              :in std_logic_vector(8 DOWNTO 0);
     Lc1189              :in std_logic_vector(8 DOWNTO 0);
     Lc1190              :in std_logic_vector(8 DOWNTO 0);
     Lc1191              :in std_logic_vector(8 DOWNTO 0);
     Lc1192              :in std_logic_vector(8 DOWNTO 0);
     Lc1193              :in std_logic_vector(8 DOWNTO 0);
     Lc1194              :in std_logic_vector(8 DOWNTO 0);
     Lc1195              :in std_logic_vector(8 DOWNTO 0);
     Lc1196              :in std_logic_vector(8 DOWNTO 0);
     Lc1197              :in std_logic_vector(8 DOWNTO 0);
     Lc1198              :in std_logic_vector(8 DOWNTO 0);
     Lc1199              :in std_logic_vector(8 DOWNTO 0);
     Lc1200              :in std_logic_vector(8 DOWNTO 0);
     Lc1201              :in std_logic_vector(8 DOWNTO 0);
     Lc1202              :in std_logic_vector(8 DOWNTO 0);
     Lc1203              :in std_logic_vector(8 DOWNTO 0);
     Lc1204              :in std_logic_vector(8 DOWNTO 0);
     Lc1205              :in std_logic_vector(8 DOWNTO 0);
     Lc1206              :in std_logic_vector(8 DOWNTO 0);
     Lc1207              :in std_logic_vector(8 DOWNTO 0);
     Lc1208              :in std_logic_vector(8 DOWNTO 0);
     Lc1209              :in std_logic_vector(8 DOWNTO 0);
     Lc1210              :in std_logic_vector(8 DOWNTO 0);
     Lc1211              :in std_logic_vector(8 DOWNTO 0);
     Lc1212              :in std_logic_vector(8 DOWNTO 0);
     Lc1213              :in std_logic_vector(8 DOWNTO 0);
     Lc1214              :in std_logic_vector(8 DOWNTO 0);
     Lc1215              :in std_logic_vector(8 DOWNTO 0);
     Lc1216              :in std_logic_vector(8 DOWNTO 0);
     Lc1217              :in std_logic_vector(8 DOWNTO 0);
     Lc1218              :in std_logic_vector(8 DOWNTO 0);
     Lc1219              :in std_logic_vector(8 DOWNTO 0);
     Lc1220              :in std_logic_vector(8 DOWNTO 0);
     Lc1221              :in std_logic_vector(8 DOWNTO 0);
     Lc1222              :in std_logic_vector(8 DOWNTO 0);
     Lc1223              :in std_logic_vector(8 DOWNTO 0);
     Lc1224              :in std_logic_vector(8 DOWNTO 0);
     Lc1225              :in std_logic_vector(8 DOWNTO 0);
     Lc1226              :in std_logic_vector(8 DOWNTO 0);
     Lc1227              :in std_logic_vector(8 DOWNTO 0);
     Lc1228              :in std_logic_vector(8 DOWNTO 0);
     Lc1229              :in std_logic_vector(8 DOWNTO 0);
     Lc1230              :in std_logic_vector(8 DOWNTO 0);
     Lc1231              :in std_logic_vector(8 DOWNTO 0);
     Lc1232              :in std_logic_vector(8 DOWNTO 0);
     Lc1233              :in std_logic_vector(8 DOWNTO 0);
     Lc1234              :in std_logic_vector(8 DOWNTO 0);
     Lc1235              :in std_logic_vector(8 DOWNTO 0);
     Lc1236              :in std_logic_vector(8 DOWNTO 0);
     Lc1237              :in std_logic_vector(8 DOWNTO 0);
     Lc1238              :in std_logic_vector(8 DOWNTO 0);
     Lc1239              :in std_logic_vector(8 DOWNTO 0);
     Lc1240              :in std_logic_vector(8 DOWNTO 0);
     Lc1241              :in std_logic_vector(8 DOWNTO 0);
     Lc1242              :in std_logic_vector(8 DOWNTO 0);
     Lc1243              :in std_logic_vector(8 DOWNTO 0);
     Lc1244              :in std_logic_vector(8 DOWNTO 0);
     Lc1245              :in std_logic_vector(8 DOWNTO 0);
     Lc1246              :in std_logic_vector(8 DOWNTO 0);
     Lc1247              :in std_logic_vector(8 DOWNTO 0);
     Lc1248              :in std_logic_vector(8 DOWNTO 0);
     Lc1249              :in std_logic_vector(8 DOWNTO 0);
     Lc1250              :in std_logic_vector(8 DOWNTO 0);
     Lc1251              :in std_logic_vector(8 DOWNTO 0);
     Lc1252              :in std_logic_vector(8 DOWNTO 0);
     Lc1253              :in std_logic_vector(8 DOWNTO 0);
     Lc1254              :in std_logic_vector(8 DOWNTO 0);
     Lc1255              :in std_logic_vector(8 DOWNTO 0);
     Lc1256              :in std_logic_vector(8 DOWNTO 0);
     Lc1257              :in std_logic_vector(8 DOWNTO 0);
     Lc1258              :in std_logic_vector(8 DOWNTO 0);
     Lc1259              :in std_logic_vector(8 DOWNTO 0);
     Lc1260              :in std_logic_vector(8 DOWNTO 0);
     Lc1261              :in std_logic_vector(8 DOWNTO 0);
     Lc1262              :in std_logic_vector(8 DOWNTO 0);
     Lc1263              :in std_logic_vector(8 DOWNTO 0);
     Lc1264              :in std_logic_vector(8 DOWNTO 0);
     Lc1265              :in std_logic_vector(8 DOWNTO 0);
     Lc1266              :in std_logic_vector(8 DOWNTO 0);
     Lc1267              :in std_logic_vector(8 DOWNTO 0);
     Lc1268              :in std_logic_vector(8 DOWNTO 0);
     Lc1269              :in std_logic_vector(8 DOWNTO 0);
     Lc1270              :in std_logic_vector(8 DOWNTO 0);
     Lc1271              :in std_logic_vector(8 DOWNTO 0);
     Lc1272              :in std_logic_vector(8 DOWNTO 0);
     Lc1273              :in std_logic_vector(8 DOWNTO 0);
     Lc1274              :in std_logic_vector(8 DOWNTO 0);
     Lc1275              :in std_logic_vector(8 DOWNTO 0);
     Lc1276              :in std_logic_vector(8 DOWNTO 0);
     Lc1277              :in std_logic_vector(8 DOWNTO 0);
     Lc1278              :in std_logic_vector(8 DOWNTO 0);
     Lc1279              :in std_logic_vector(8 DOWNTO 0);
     Lc1280              :in std_logic_vector(8 DOWNTO 0);
     Lc1281              :in std_logic_vector(8 DOWNTO 0);
     Lc1282              :in std_logic_vector(8 DOWNTO 0);
     Lc1283              :in std_logic_vector(8 DOWNTO 0);
     Lc1284              :in std_logic_vector(8 DOWNTO 0);
     Lc1285              :in std_logic_vector(8 DOWNTO 0);
     Lc1286              :in std_logic_vector(8 DOWNTO 0);
     Lc1287              :in std_logic_vector(8 DOWNTO 0);
     Lc1288              :in std_logic_vector(8 DOWNTO 0);
     Lc1289              :in std_logic_vector(8 DOWNTO 0);
     Lc1290              :in std_logic_vector(8 DOWNTO 0);
     Lc1291              :in std_logic_vector(8 DOWNTO 0);
     Lc1292              :in std_logic_vector(8 DOWNTO 0);
     Lc1293              :in std_logic_vector(8 DOWNTO 0);
     Lc1294              :in std_logic_vector(8 DOWNTO 0);
     Lc1295              :in std_logic_vector(8 DOWNTO 0);
     Lc1296              :in std_logic_vector(8 DOWNTO 0);
     Lc1297              :in std_logic_vector(8 DOWNTO 0);
     Lc1298              :in std_logic_vector(8 DOWNTO 0);
     Lc1299              :in std_logic_vector(8 DOWNTO 0);
     Lc1300              :in std_logic_vector(8 DOWNTO 0);
     Lc1301              :in std_logic_vector(8 DOWNTO 0);
     Lc1302              :in std_logic_vector(8 DOWNTO 0);
     Lc1303              :in std_logic_vector(8 DOWNTO 0);
     Lc1304              :in std_logic_vector(8 DOWNTO 0);
     Lc1305              :in std_logic_vector(8 DOWNTO 0);
     Lc1306              :in std_logic_vector(8 DOWNTO 0);
     Lc1307              :in std_logic_vector(8 DOWNTO 0);
     Lc1308              :in std_logic_vector(8 DOWNTO 0);
     Lc1309              :in std_logic_vector(8 DOWNTO 0);
     Lc1310              :in std_logic_vector(8 DOWNTO 0);
     Lc1311              :in std_logic_vector(8 DOWNTO 0);
     Lc1312              :in std_logic_vector(8 DOWNTO 0);
     Lc1313              :in std_logic_vector(8 DOWNTO 0);
     Lc1314              :in std_logic_vector(8 DOWNTO 0);
     Lc1315              :in std_logic_vector(8 DOWNTO 0);
     Lc1316              :in std_logic_vector(8 DOWNTO 0);
     Lc1317              :in std_logic_vector(8 DOWNTO 0);
     Lc1318              :in std_logic_vector(8 DOWNTO 0);
     Lc1319              :in std_logic_vector(8 DOWNTO 0);
     Lc1320              :in std_logic_vector(8 DOWNTO 0);
     Lc1321              :in std_logic_vector(8 DOWNTO 0);
     Lc1322              :in std_logic_vector(8 DOWNTO 0);
     Lc1323              :in std_logic_vector(8 DOWNTO 0);
     Lc1324              :in std_logic_vector(8 DOWNTO 0);
     Lc1325              :in std_logic_vector(8 DOWNTO 0);
     Lc1326              :in std_logic_vector(8 DOWNTO 0);
     Lc1327              :in std_logic_vector(8 DOWNTO 0);
     Lc1328              :in std_logic_vector(8 DOWNTO 0);
     Lc1329              :in std_logic_vector(8 DOWNTO 0);
     Lc1330              :in std_logic_vector(8 DOWNTO 0);
     Lc1331              :in std_logic_vector(8 DOWNTO 0);
     Lc1332              :in std_logic_vector(8 DOWNTO 0);
     Lc1333              :in std_logic_vector(8 DOWNTO 0);
     Lc1334              :in std_logic_vector(8 DOWNTO 0);
     Lc1335              :in std_logic_vector(8 DOWNTO 0);
     Lc1336              :in std_logic_vector(8 DOWNTO 0);
     Lc1337              :in std_logic_vector(8 DOWNTO 0);
     Lc1338              :in std_logic_vector(8 DOWNTO 0);
     Lc1339              :in std_logic_vector(8 DOWNTO 0);
     Lc1340              :in std_logic_vector(8 DOWNTO 0);
     Lc1341              :in std_logic_vector(8 DOWNTO 0);
     Lc1342              :in std_logic_vector(8 DOWNTO 0);
     Lc1343              :in std_logic_vector(8 DOWNTO 0);
     Lc1344              :in std_logic_vector(8 DOWNTO 0);
     Lc1345              :in std_logic_vector(8 DOWNTO 0);
     Lc1346              :in std_logic_vector(8 DOWNTO 0);
     Lc1347              :in std_logic_vector(8 DOWNTO 0);
     Lc1348              :in std_logic_vector(8 DOWNTO 0);
     Lc1349              :in std_logic_vector(8 DOWNTO 0);
     Lc1350              :in std_logic_vector(8 DOWNTO 0);
     Lc1351              :in std_logic_vector(8 DOWNTO 0);
     Lc1352              :in std_logic_vector(8 DOWNTO 0);
     Lc1353              :in std_logic_vector(8 DOWNTO 0);
     Lc1354              :in std_logic_vector(8 DOWNTO 0);
     Lc1355              :in std_logic_vector(8 DOWNTO 0);
     Lc1356              :in std_logic_vector(8 DOWNTO 0);
     Lc1357              :in std_logic_vector(8 DOWNTO 0);
     Lc1358              :in std_logic_vector(8 DOWNTO 0);
     Lc1359              :in std_logic_vector(8 DOWNTO 0);
     Lc1360              :in std_logic_vector(8 DOWNTO 0);
     Lc1361              :in std_logic_vector(8 DOWNTO 0);
     Lc1362              :in std_logic_vector(8 DOWNTO 0);
     Lc1363              :in std_logic_vector(8 DOWNTO 0);
     Lc1364              :in std_logic_vector(8 DOWNTO 0);
     Lc1365              :in std_logic_vector(8 DOWNTO 0);
     Lc1366              :in std_logic_vector(8 DOWNTO 0);
     Lc1367              :in std_logic_vector(8 DOWNTO 0);
     Lc1368              :in std_logic_vector(8 DOWNTO 0);
     Lc1369              :in std_logic_vector(8 DOWNTO 0);
     Lc1370              :in std_logic_vector(8 DOWNTO 0);
     Lc1371              :in std_logic_vector(8 DOWNTO 0);
     Lc1372              :in std_logic_vector(8 DOWNTO 0);
     Lc1373              :in std_logic_vector(8 DOWNTO 0);
     Lc1374              :in std_logic_vector(8 DOWNTO 0);
     Lc1375              :in std_logic_vector(8 DOWNTO 0);
     Lc1376              :in std_logic_vector(8 DOWNTO 0);
     Lc1377              :in std_logic_vector(8 DOWNTO 0);
     Lc1378              :in std_logic_vector(8 DOWNTO 0);
     Lc1379              :in std_logic_vector(8 DOWNTO 0);
     Lc1380              :in std_logic_vector(8 DOWNTO 0);
     Lc1381              :in std_logic_vector(8 DOWNTO 0);
     Lc1382              :in std_logic_vector(8 DOWNTO 0);
     Lc1383              :in std_logic_vector(8 DOWNTO 0);
     Lc1384              :in std_logic_vector(8 DOWNTO 0);
     Lc1385              :in std_logic_vector(8 DOWNTO 0);
     Lc1386              :in std_logic_vector(8 DOWNTO 0);
     Lc1387              :in std_logic_vector(8 DOWNTO 0);
     Lc1388              :in std_logic_vector(8 DOWNTO 0);
     Lc1389              :in std_logic_vector(8 DOWNTO 0);
     Lc1390              :in std_logic_vector(8 DOWNTO 0);
     Lc1391              :in std_logic_vector(8 DOWNTO 0);
     Lc1392              :in std_logic_vector(8 DOWNTO 0);
     Lc1393              :in std_logic_vector(8 DOWNTO 0);
     Lc1394              :in std_logic_vector(8 DOWNTO 0);
     Lc1395              :in std_logic_vector(8 DOWNTO 0);
     Lc1396              :in std_logic_vector(8 DOWNTO 0);
     Lc1397              :in std_logic_vector(8 DOWNTO 0);
     Lc1398              :in std_logic_vector(8 DOWNTO 0);
     Lc1399              :in std_logic_vector(8 DOWNTO 0);
     Lc1400              :in std_logic_vector(8 DOWNTO 0);
     Lc1401              :in std_logic_vector(8 DOWNTO 0);
     Lc1402              :in std_logic_vector(8 DOWNTO 0);
     Lc1403              :in std_logic_vector(8 DOWNTO 0);
     Lc1404              :in std_logic_vector(8 DOWNTO 0);
     Lc1405              :in std_logic_vector(8 DOWNTO 0);
     Lc1406              :in std_logic_vector(8 DOWNTO 0);
     Lc1407              :in std_logic_vector(8 DOWNTO 0);
     Lc1408              :in std_logic_vector(8 DOWNTO 0);
     Lc1409              :in std_logic_vector(8 DOWNTO 0);
     Lc1410              :in std_logic_vector(8 DOWNTO 0);
     Lc1411              :in std_logic_vector(8 DOWNTO 0);
     Lc1412              :in std_logic_vector(8 DOWNTO 0);
     Lc1413              :in std_logic_vector(8 DOWNTO 0);
     Lc1414              :in std_logic_vector(8 DOWNTO 0);
     Lc1415              :in std_logic_vector(8 DOWNTO 0);
     Lc1416              :in std_logic_vector(8 DOWNTO 0);
     Lc1417              :in std_logic_vector(8 DOWNTO 0);
     Lc1418              :in std_logic_vector(8 DOWNTO 0);
     Lc1419              :in std_logic_vector(8 DOWNTO 0);
     Lc1420              :in std_logic_vector(8 DOWNTO 0);
     Lc1421              :in std_logic_vector(8 DOWNTO 0);
     Lc1422              :in std_logic_vector(8 DOWNTO 0);
     Lc1423              :in std_logic_vector(8 DOWNTO 0);
     Lc1424              :in std_logic_vector(8 DOWNTO 0);
     Lc1425              :in std_logic_vector(8 DOWNTO 0);
     Lc1426              :in std_logic_vector(8 DOWNTO 0);
     Lc1427              :in std_logic_vector(8 DOWNTO 0);
     Lc1428              :in std_logic_vector(8 DOWNTO 0);
     Lc1429              :in std_logic_vector(8 DOWNTO 0);
     Lc1430              :in std_logic_vector(8 DOWNTO 0);
     Lc1431              :in std_logic_vector(8 DOWNTO 0);
     Lc1432              :in std_logic_vector(8 DOWNTO 0);
     Lc1433              :in std_logic_vector(8 DOWNTO 0);
     Lc1434              :in std_logic_vector(8 DOWNTO 0);
     Lc1435              :in std_logic_vector(8 DOWNTO 0);
     Lc1436              :in std_logic_vector(8 DOWNTO 0);
     Lc1437              :in std_logic_vector(8 DOWNTO 0);
     Lc1438              :in std_logic_vector(8 DOWNTO 0);
     Lc1439              :in std_logic_vector(8 DOWNTO 0);
     Lc1440              :in std_logic_vector(8 DOWNTO 0);
     Lc1441              :in std_logic_vector(8 DOWNTO 0);
     Lc1442              :in std_logic_vector(8 DOWNTO 0);
     Lc1443              :in std_logic_vector(8 DOWNTO 0);
     Lc1444              :in std_logic_vector(8 DOWNTO 0);
     Lc1445              :in std_logic_vector(8 DOWNTO 0);
     Lc1446              :in std_logic_vector(8 DOWNTO 0);
     Lc1447              :in std_logic_vector(8 DOWNTO 0);
     Lc1448              :in std_logic_vector(8 DOWNTO 0);
     Lc1449              :in std_logic_vector(8 DOWNTO 0);
     Lc1450              :in std_logic_vector(8 DOWNTO 0);
     Lc1451              :in std_logic_vector(8 DOWNTO 0);
     Lc1452              :in std_logic_vector(8 DOWNTO 0);
     Lc1453              :in std_logic_vector(8 DOWNTO 0);
     Lc1454              :in std_logic_vector(8 DOWNTO 0);
     Lc1455              :in std_logic_vector(8 DOWNTO 0);
     Lc1456              :in std_logic_vector(8 DOWNTO 0);
     Lc1457              :in std_logic_vector(8 DOWNTO 0);
     Lc1458              :in std_logic_vector(8 DOWNTO 0);
     Lc1459              :in std_logic_vector(8 DOWNTO 0);
     Lc1460              :in std_logic_vector(8 DOWNTO 0);
     Lc1461              :in std_logic_vector(8 DOWNTO 0);
     Lc1462              :in std_logic_vector(8 DOWNTO 0);
     Lc1463              :in std_logic_vector(8 DOWNTO 0);
     Lc1464              :in std_logic_vector(8 DOWNTO 0);
     Lc1465              :in std_logic_vector(8 DOWNTO 0);
     Lc1466              :in std_logic_vector(8 DOWNTO 0);
     Lc1467              :in std_logic_vector(8 DOWNTO 0);
     Lc1468              :in std_logic_vector(8 DOWNTO 0);
     Lc1469              :in std_logic_vector(8 DOWNTO 0);
     Lc1470              :in std_logic_vector(8 DOWNTO 0);
     Lc1471              :in std_logic_vector(8 DOWNTO 0);
     Lc1472              :in std_logic_vector(8 DOWNTO 0);
     Lc1473              :in std_logic_vector(8 DOWNTO 0);
     Lc1474              :in std_logic_vector(8 DOWNTO 0);
     Lc1475              :in std_logic_vector(8 DOWNTO 0);
     Lc1476              :in std_logic_vector(8 DOWNTO 0);
     Lc1477              :in std_logic_vector(8 DOWNTO 0);
     Lc1478              :in std_logic_vector(8 DOWNTO 0);
     Lc1479              :in std_logic_vector(8 DOWNTO 0);
     Lc1480              :in std_logic_vector(8 DOWNTO 0);
     Lc1481              :in std_logic_vector(8 DOWNTO 0);
     Lc1482              :in std_logic_vector(8 DOWNTO 0);
     Lc1483              :in std_logic_vector(8 DOWNTO 0);
     Lc1484              :in std_logic_vector(8 DOWNTO 0);
     Lc1485              :in std_logic_vector(8 DOWNTO 0);
     Lc1486              :in std_logic_vector(8 DOWNTO 0);
     Lc1487              :in std_logic_vector(8 DOWNTO 0);
     Lc1488              :in std_logic_vector(8 DOWNTO 0);
     Lc1489              :in std_logic_vector(8 DOWNTO 0);
     Lc1490              :in std_logic_vector(8 DOWNTO 0);
     Lc1491              :in std_logic_vector(8 DOWNTO 0);
     Lc1492              :in std_logic_vector(8 DOWNTO 0);
     Lc1493              :in std_logic_vector(8 DOWNTO 0);
     Lc1494              :in std_logic_vector(8 DOWNTO 0);
     Lc1495              :in std_logic_vector(8 DOWNTO 0);
     Lc1496              :in std_logic_vector(8 DOWNTO 0);
     Lc1497              :in std_logic_vector(8 DOWNTO 0);
     Lc1498              :in std_logic_vector(8 DOWNTO 0);
     Lc1499              :in std_logic_vector(8 DOWNTO 0);
     Lc1500              :in std_logic_vector(8 DOWNTO 0);
     Lc1501              :in std_logic_vector(8 DOWNTO 0);
     Lc1502              :in std_logic_vector(8 DOWNTO 0);
     Lc1503              :in std_logic_vector(8 DOWNTO 0);
     Lc1504              :in std_logic_vector(8 DOWNTO 0);
     Lc1505              :in std_logic_vector(8 DOWNTO 0);
     Lc1506              :in std_logic_vector(8 DOWNTO 0);
     Lc1507              :in std_logic_vector(8 DOWNTO 0);
     Lc1508              :in std_logic_vector(8 DOWNTO 0);
     Lc1509              :in std_logic_vector(8 DOWNTO 0);
     Lc1510              :in std_logic_vector(8 DOWNTO 0);
     Lc1511              :in std_logic_vector(8 DOWNTO 0);
     Lc1512              :in std_logic_vector(8 DOWNTO 0);
     Lc1513              :in std_logic_vector(8 DOWNTO 0);
     Lc1514              :in std_logic_vector(8 DOWNTO 0);
     Lc1515              :in std_logic_vector(8 DOWNTO 0);
     Lc1516              :in std_logic_vector(8 DOWNTO 0);
     Lc1517              :in std_logic_vector(8 DOWNTO 0);
     Lc1518              :in std_logic_vector(8 DOWNTO 0);
     Lc1519              :in std_logic_vector(8 DOWNTO 0);
     Lc1520              :in std_logic_vector(8 DOWNTO 0);
     Lc1521              :in std_logic_vector(8 DOWNTO 0);
     Lc1522              :in std_logic_vector(8 DOWNTO 0);
     Lc1523              :in std_logic_vector(8 DOWNTO 0);
     Lc1524              :in std_logic_vector(8 DOWNTO 0);
     Lc1525              :in std_logic_vector(8 DOWNTO 0);
     Lc1526              :in std_logic_vector(8 DOWNTO 0);
     Lc1527              :in std_logic_vector(8 DOWNTO 0);
     Lc1528              :in std_logic_vector(8 DOWNTO 0);
     Lc1529              :in std_logic_vector(8 DOWNTO 0);
     Lc1530              :in std_logic_vector(8 DOWNTO 0);
     Lc1531              :in std_logic_vector(8 DOWNTO 0);
     Lc1532              :in std_logic_vector(8 DOWNTO 0);
     Lc1533              :in std_logic_vector(8 DOWNTO 0);
     Lc1534              :in std_logic_vector(8 DOWNTO 0);
     Lc1535              :in std_logic_vector(8 DOWNTO 0);
     Lc1536              :in std_logic_vector(8 DOWNTO 0);
     Lc1537              :in std_logic_vector(8 DOWNTO 0);
     Lc1538              :in std_logic_vector(8 DOWNTO 0);
     Lc1539              :in std_logic_vector(8 DOWNTO 0);
     Lc1540              :in std_logic_vector(8 DOWNTO 0);
     Lc1541              :in std_logic_vector(8 DOWNTO 0);
     Lc1542              :in std_logic_vector(8 DOWNTO 0);
     Lc1543              :in std_logic_vector(8 DOWNTO 0);
     Lc1544              :in std_logic_vector(8 DOWNTO 0);
     Lc1545              :in std_logic_vector(8 DOWNTO 0);
     Lc1546              :in std_logic_vector(8 DOWNTO 0);
     Lc1547              :in std_logic_vector(8 DOWNTO 0);
     Lc1548              :in std_logic_vector(8 DOWNTO 0);
     Lc1549              :in std_logic_vector(8 DOWNTO 0);
     Lc1550              :in std_logic_vector(8 DOWNTO 0);
     Lc1551              :in std_logic_vector(8 DOWNTO 0);
     Lc1552              :in std_logic_vector(8 DOWNTO 0);
     Lc1553              :in std_logic_vector(8 DOWNTO 0);
     Lc1554              :in std_logic_vector(8 DOWNTO 0);
     Lc1555              :in std_logic_vector(8 DOWNTO 0);
     Lc1556              :in std_logic_vector(8 DOWNTO 0);
     Lc1557              :in std_logic_vector(8 DOWNTO 0);
     Lc1558              :in std_logic_vector(8 DOWNTO 0);
     Lc1559              :in std_logic_vector(8 DOWNTO 0);
     Lc1560              :in std_logic_vector(8 DOWNTO 0);
     Lc1561              :in std_logic_vector(8 DOWNTO 0);
     Lc1562              :in std_logic_vector(8 DOWNTO 0);
     Lc1563              :in std_logic_vector(8 DOWNTO 0);
     Lc1564              :in std_logic_vector(8 DOWNTO 0);
     Lc1565              :in std_logic_vector(8 DOWNTO 0);
     Lc1566              :in std_logic_vector(8 DOWNTO 0);
     Lc1567              :in std_logic_vector(8 DOWNTO 0);
     Lc1568              :in std_logic_vector(8 DOWNTO 0);
     Lc1569              :in std_logic_vector(8 DOWNTO 0);
     Lc1570              :in std_logic_vector(8 DOWNTO 0);
     Lc1571              :in std_logic_vector(8 DOWNTO 0);
     Lc1572              :in std_logic_vector(8 DOWNTO 0);
     Lc1573              :in std_logic_vector(8 DOWNTO 0);
     Lc1574              :in std_logic_vector(8 DOWNTO 0);
     Lc1575              :in std_logic_vector(8 DOWNTO 0);
     Lc1576              :in std_logic_vector(8 DOWNTO 0);
     Lc1577              :in std_logic_vector(8 DOWNTO 0);
     Lc1578              :in std_logic_vector(8 DOWNTO 0);
     Lc1579              :in std_logic_vector(8 DOWNTO 0);
     Lc1580              :in std_logic_vector(8 DOWNTO 0);
     Lc1581              :in std_logic_vector(8 DOWNTO 0);
     Lc1582              :in std_logic_vector(8 DOWNTO 0);
     Lc1583              :in std_logic_vector(8 DOWNTO 0);
     Lc1584              :in std_logic_vector(8 DOWNTO 0);
     Lc1585              :in std_logic_vector(8 DOWNTO 0);
     Lc1586              :in std_logic_vector(8 DOWNTO 0);
     Lc1587              :in std_logic_vector(8 DOWNTO 0);
     Lc1588              :in std_logic_vector(8 DOWNTO 0);
     Lc1589              :in std_logic_vector(8 DOWNTO 0);
     Lc1590              :in std_logic_vector(8 DOWNTO 0);
     Lc1591              :in std_logic_vector(8 DOWNTO 0);
     Lc1592              :in std_logic_vector(8 DOWNTO 0);
     Lc1593              :in std_logic_vector(8 DOWNTO 0);
     Lc1594              :in std_logic_vector(8 DOWNTO 0);
     Lc1595              :in std_logic_vector(8 DOWNTO 0);
     Lc1596              :in std_logic_vector(8 DOWNTO 0);
     Lc1597              :in std_logic_vector(8 DOWNTO 0);
     Lc1598              :in std_logic_vector(8 DOWNTO 0);
     Lc1599              :in std_logic_vector(8 DOWNTO 0);
     Lc1600              :in std_logic_vector(8 DOWNTO 0);
     Lc1601              :in std_logic_vector(8 DOWNTO 0);
     Lc1602              :in std_logic_vector(8 DOWNTO 0);
     Lc1603              :in std_logic_vector(8 DOWNTO 0);
     Lc1604              :in std_logic_vector(8 DOWNTO 0);
     Lc1605              :in std_logic_vector(8 DOWNTO 0);
     Lc1606              :in std_logic_vector(8 DOWNTO 0);
     Lc1607              :in std_logic_vector(8 DOWNTO 0);
     Lc1608              :in std_logic_vector(8 DOWNTO 0);
     Lc1609              :in std_logic_vector(8 DOWNTO 0);
     Lc1610              :in std_logic_vector(8 DOWNTO 0);
     Lc1611              :in std_logic_vector(8 DOWNTO 0);
     Lc1612              :in std_logic_vector(8 DOWNTO 0);
     Lc1613              :in std_logic_vector(8 DOWNTO 0);
     Lc1614              :in std_logic_vector(8 DOWNTO 0);
     Lc1615              :in std_logic_vector(8 DOWNTO 0);
     Lc1616              :in std_logic_vector(8 DOWNTO 0);
     Lc1617              :in std_logic_vector(8 DOWNTO 0);
     Lc1618              :in std_logic_vector(8 DOWNTO 0);
     Lc1619              :in std_logic_vector(8 DOWNTO 0);
     Lc1620              :in std_logic_vector(8 DOWNTO 0);
     Lc1621              :in std_logic_vector(8 DOWNTO 0);
     Lc1622              :in std_logic_vector(8 DOWNTO 0);
     Lc1623              :in std_logic_vector(8 DOWNTO 0);
     Lc1624              :in std_logic_vector(8 DOWNTO 0);
     Lc1625              :in std_logic_vector(8 DOWNTO 0);
     Lc1626              :in std_logic_vector(8 DOWNTO 0);
     Lc1627              :in std_logic_vector(8 DOWNTO 0);
     Lc1628              :in std_logic_vector(8 DOWNTO 0);
     Lc1629              :in std_logic_vector(8 DOWNTO 0);
     Lc1630              :in std_logic_vector(8 DOWNTO 0);
     Lc1631              :in std_logic_vector(8 DOWNTO 0);
     Lc1632              :in std_logic_vector(8 DOWNTO 0);
     Lc1633              :in std_logic_vector(8 DOWNTO 0);
     Lc1634              :in std_logic_vector(8 DOWNTO 0);
     Lc1635              :in std_logic_vector(8 DOWNTO 0);
     Lc1636              :in std_logic_vector(8 DOWNTO 0);
     Lc1637              :in std_logic_vector(8 DOWNTO 0);
     Lc1638              :in std_logic_vector(8 DOWNTO 0);
     Lc1639              :in std_logic_vector(8 DOWNTO 0);
     Lc1640              :in std_logic_vector(8 DOWNTO 0);
     Lc1641              :in std_logic_vector(8 DOWNTO 0);
     Lc1642              :in std_logic_vector(8 DOWNTO 0);
     Lc1643              :in std_logic_vector(8 DOWNTO 0);
     Lc1644              :in std_logic_vector(8 DOWNTO 0);
     Lc1645              :in std_logic_vector(8 DOWNTO 0);
     Lc1646              :in std_logic_vector(8 DOWNTO 0);
     Lc1647              :in std_logic_vector(8 DOWNTO 0);
     Lc1648              :in std_logic_vector(8 DOWNTO 0);
     Lc1649              :in std_logic_vector(8 DOWNTO 0);
     Lc1650              :in std_logic_vector(8 DOWNTO 0);
     Lc1651              :in std_logic_vector(8 DOWNTO 0);
     Lc1652              :in std_logic_vector(8 DOWNTO 0);
     Lc1653              :in std_logic_vector(8 DOWNTO 0);
     Lc1654              :in std_logic_vector(8 DOWNTO 0);
     Lc1655              :in std_logic_vector(8 DOWNTO 0);
     Lc1656              :in std_logic_vector(8 DOWNTO 0);
     Lc1657              :in std_logic_vector(8 DOWNTO 0);
     Lc1658              :in std_logic_vector(8 DOWNTO 0);
     Lc1659              :in std_logic_vector(8 DOWNTO 0);
     Lc1660              :in std_logic_vector(8 DOWNTO 0);
     Lc1661              :in std_logic_vector(8 DOWNTO 0);
     Lc1662              :in std_logic_vector(8 DOWNTO 0);
     Lc1663              :in std_logic_vector(8 DOWNTO 0);
     Lc1664              :in std_logic_vector(8 DOWNTO 0);
     Lc1665              :in std_logic_vector(8 DOWNTO 0);
     Lc1666              :in std_logic_vector(8 DOWNTO 0);
     Lc1667              :in std_logic_vector(8 DOWNTO 0);
     Lc1668              :in std_logic_vector(8 DOWNTO 0);
     Lc1669              :in std_logic_vector(8 DOWNTO 0);
     Lc1670              :in std_logic_vector(8 DOWNTO 0);
     Lc1671              :in std_logic_vector(8 DOWNTO 0);
     Lc1672              :in std_logic_vector(8 DOWNTO 0);
     Lc1673              :in std_logic_vector(8 DOWNTO 0);
     Lc1674              :in std_logic_vector(8 DOWNTO 0);
     Lc1675              :in std_logic_vector(8 DOWNTO 0);
     Lc1676              :in std_logic_vector(8 DOWNTO 0);
     Lc1677              :in std_logic_vector(8 DOWNTO 0);
     Lc1678              :in std_logic_vector(8 DOWNTO 0);
     Lc1679              :in std_logic_vector(8 DOWNTO 0);
     Lc1680              :in std_logic_vector(8 DOWNTO 0);
     Lc1681              :in std_logic_vector(8 DOWNTO 0);
     Lc1682              :in std_logic_vector(8 DOWNTO 0);
     Lc1683              :in std_logic_vector(8 DOWNTO 0);
     Lc1684              :in std_logic_vector(8 DOWNTO 0);
     Lc1685              :in std_logic_vector(8 DOWNTO 0);
     Lc1686              :in std_logic_vector(8 DOWNTO 0);
     Lc1687              :in std_logic_vector(8 DOWNTO 0);
     Lc1688              :in std_logic_vector(8 DOWNTO 0);
     Lc1689              :in std_logic_vector(8 DOWNTO 0);
     Lc1690              :in std_logic_vector(8 DOWNTO 0);
     Lc1691              :in std_logic_vector(8 DOWNTO 0);
     Lc1692              :in std_logic_vector(8 DOWNTO 0);
     Lc1693              :in std_logic_vector(8 DOWNTO 0);
     Lc1694              :in std_logic_vector(8 DOWNTO 0);
     Lc1695              :in std_logic_vector(8 DOWNTO 0);
     Lc1696              :in std_logic_vector(8 DOWNTO 0);
     Lc1697              :in std_logic_vector(8 DOWNTO 0);
     Lc1698              :in std_logic_vector(8 DOWNTO 0);
     Lc1699              :in std_logic_vector(8 DOWNTO 0);
     Lc1700              :in std_logic_vector(8 DOWNTO 0);
     Lc1701              :in std_logic_vector(8 DOWNTO 0);
     Lc1702              :in std_logic_vector(8 DOWNTO 0);
     Lc1703              :in std_logic_vector(8 DOWNTO 0);
     Lc1704              :in std_logic_vector(8 DOWNTO 0);
     Lc1705              :in std_logic_vector(8 DOWNTO 0);
     Lc1706              :in std_logic_vector(8 DOWNTO 0);
     Lc1707              :in std_logic_vector(8 DOWNTO 0);
     Lc1708              :in std_logic_vector(8 DOWNTO 0);
     Lc1709              :in std_logic_vector(8 DOWNTO 0);
     Lc1710              :in std_logic_vector(8 DOWNTO 0);
     Lc1711              :in std_logic_vector(8 DOWNTO 0);
     Lc1712              :in std_logic_vector(8 DOWNTO 0);
     Lc1713              :in std_logic_vector(8 DOWNTO 0);
     Lc1714              :in std_logic_vector(8 DOWNTO 0);
     Lc1715              :in std_logic_vector(8 DOWNTO 0);
     Lc1716              :in std_logic_vector(8 DOWNTO 0);
     Lc1717              :in std_logic_vector(8 DOWNTO 0);
     Lc1718              :in std_logic_vector(8 DOWNTO 0);
     Lc1719              :in std_logic_vector(8 DOWNTO 0);
     Lc1720              :in std_logic_vector(8 DOWNTO 0);
     Lc1721              :in std_logic_vector(8 DOWNTO 0);
     Lc1722              :in std_logic_vector(8 DOWNTO 0);
     Lc1723              :in std_logic_vector(8 DOWNTO 0);
     Lc1724              :in std_logic_vector(8 DOWNTO 0);
     Lc1725              :in std_logic_vector(8 DOWNTO 0);
     Lc1726              :in std_logic_vector(8 DOWNTO 0);
     Lc1727              :in std_logic_vector(8 DOWNTO 0);
     Lc1728              :in std_logic_vector(8 DOWNTO 0);
     Lc1729              :in std_logic_vector(8 DOWNTO 0);
     Lc1730              :in std_logic_vector(8 DOWNTO 0);
     Lc1731              :in std_logic_vector(8 DOWNTO 0);
     Lc1732              :in std_logic_vector(8 DOWNTO 0);
     Lc1733              :in std_logic_vector(8 DOWNTO 0);
     Lc1734              :in std_logic_vector(8 DOWNTO 0);
     Lc1735              :in std_logic_vector(8 DOWNTO 0);
     Lc1736              :in std_logic_vector(8 DOWNTO 0);
     Lc1737              :in std_logic_vector(8 DOWNTO 0);
     Lc1738              :in std_logic_vector(8 DOWNTO 0);
     Lc1739              :in std_logic_vector(8 DOWNTO 0);
     Lc1740              :in std_logic_vector(8 DOWNTO 0);
     Lc1741              :in std_logic_vector(8 DOWNTO 0);
     Lc1742              :in std_logic_vector(8 DOWNTO 0);
     Lc1743              :in std_logic_vector(8 DOWNTO 0);
     Lc1744              :in std_logic_vector(8 DOWNTO 0);
     Lc1745              :in std_logic_vector(8 DOWNTO 0);
     Lc1746              :in std_logic_vector(8 DOWNTO 0);
     Lc1747              :in std_logic_vector(8 DOWNTO 0);
     Lc1748              :in std_logic_vector(8 DOWNTO 0);
     Lc1749              :in std_logic_vector(8 DOWNTO 0);
     Lc1750              :in std_logic_vector(8 DOWNTO 0);
     Lc1751              :in std_logic_vector(8 DOWNTO 0);
     Lc1752              :in std_logic_vector(8 DOWNTO 0);
     Lc1753              :in std_logic_vector(8 DOWNTO 0);
     Lc1754              :in std_logic_vector(8 DOWNTO 0);
     Lc1755              :in std_logic_vector(8 DOWNTO 0);
     Lc1756              :in std_logic_vector(8 DOWNTO 0);
     Lc1757              :in std_logic_vector(8 DOWNTO 0);
     Lc1758              :in std_logic_vector(8 DOWNTO 0);
     Lc1759              :in std_logic_vector(8 DOWNTO 0);
     Lc1760              :in std_logic_vector(8 DOWNTO 0);
     Lc1761              :in std_logic_vector(8 DOWNTO 0);
     Lc1762              :in std_logic_vector(8 DOWNTO 0);
     Lc1763              :in std_logic_vector(8 DOWNTO 0);
     Lc1764              :in std_logic_vector(8 DOWNTO 0);
     Lc1765              :in std_logic_vector(8 DOWNTO 0);
     Lc1766              :in std_logic_vector(8 DOWNTO 0);
     Lc1767              :in std_logic_vector(8 DOWNTO 0);
     Lc1768              :in std_logic_vector(8 DOWNTO 0);
     Lc1769              :in std_logic_vector(8 DOWNTO 0);
     Lc1770              :in std_logic_vector(8 DOWNTO 0);
     Lc1771              :in std_logic_vector(8 DOWNTO 0);
     Lc1772              :in std_logic_vector(8 DOWNTO 0);
     Lc1773              :in std_logic_vector(8 DOWNTO 0);
     Lc1774              :in std_logic_vector(8 DOWNTO 0);
     Lc1775              :in std_logic_vector(8 DOWNTO 0);
     Lc1776              :in std_logic_vector(8 DOWNTO 0);
     Lc1777              :in std_logic_vector(8 DOWNTO 0);
     Lc1778              :in std_logic_vector(8 DOWNTO 0);
     Lc1779              :in std_logic_vector(8 DOWNTO 0);
     Lc1780              :in std_logic_vector(8 DOWNTO 0);
     Lc1781              :in std_logic_vector(8 DOWNTO 0);
     Lc1782              :in std_logic_vector(8 DOWNTO 0);
     Lc1783              :in std_logic_vector(8 DOWNTO 0);
     Lc1784              :in std_logic_vector(8 DOWNTO 0);
     Lc1785              :in std_logic_vector(8 DOWNTO 0);
     Lc1786              :in std_logic_vector(8 DOWNTO 0);
     Lc1787              :in std_logic_vector(8 DOWNTO 0);
     Lc1788              :in std_logic_vector(8 DOWNTO 0);
     Lc1789              :in std_logic_vector(8 DOWNTO 0);
     Lc1790              :in std_logic_vector(8 DOWNTO 0);
     Lc1791              :in std_logic_vector(8 DOWNTO 0);
     Lc1792              :in std_logic_vector(8 DOWNTO 0);
     Lc1793              :in std_logic_vector(8 DOWNTO 0);
     Lc1794              :in std_logic_vector(8 DOWNTO 0);
     Lc1795              :in std_logic_vector(8 DOWNTO 0);
     Lc1796              :in std_logic_vector(8 DOWNTO 0);
     Lc1797              :in std_logic_vector(8 DOWNTO 0);
     Lc1798              :in std_logic_vector(8 DOWNTO 0);
     Lc1799              :in std_logic_vector(8 DOWNTO 0);
     Lc1800              :in std_logic_vector(8 DOWNTO 0);
     Lc1801              :in std_logic_vector(8 DOWNTO 0);
     Lc1802              :in std_logic_vector(8 DOWNTO 0);
     Lc1803              :in std_logic_vector(8 DOWNTO 0);
     Lc1804              :in std_logic_vector(8 DOWNTO 0);
     Lc1805              :in std_logic_vector(8 DOWNTO 0);
     Lc1806              :in std_logic_vector(8 DOWNTO 0);
     Lc1807              :in std_logic_vector(8 DOWNTO 0);
     Lc1808              :in std_logic_vector(8 DOWNTO 0);
     Lc1809              :in std_logic_vector(8 DOWNTO 0);
     Lc1810              :in std_logic_vector(8 DOWNTO 0);
     Lc1811              :in std_logic_vector(8 DOWNTO 0);
     Lc1812              :in std_logic_vector(8 DOWNTO 0);
     Lc1813              :in std_logic_vector(8 DOWNTO 0);
     Lc1814              :in std_logic_vector(8 DOWNTO 0);
     Lc1815              :in std_logic_vector(8 DOWNTO 0);
     Lc1816              :in std_logic_vector(8 DOWNTO 0);
     Lc1817              :in std_logic_vector(8 DOWNTO 0);
     Lc1818              :in std_logic_vector(8 DOWNTO 0);
     Lc1819              :in std_logic_vector(8 DOWNTO 0);
     Lc1820              :in std_logic_vector(8 DOWNTO 0);
     Lc1821              :in std_logic_vector(8 DOWNTO 0);
     Lc1822              :in std_logic_vector(8 DOWNTO 0);
     Lc1823              :in std_logic_vector(8 DOWNTO 0);
     Lc1824              :in std_logic_vector(8 DOWNTO 0);
     Lc1825              :in std_logic_vector(8 DOWNTO 0);
     Lc1826              :in std_logic_vector(8 DOWNTO 0);
     Lc1827              :in std_logic_vector(8 DOWNTO 0);
     Lc1828              :in std_logic_vector(8 DOWNTO 0);
     Lc1829              :in std_logic_vector(8 DOWNTO 0);
     Lc1830              :in std_logic_vector(8 DOWNTO 0);
     Lc1831              :in std_logic_vector(8 DOWNTO 0);
     Lc1832              :in std_logic_vector(8 DOWNTO 0);
     Lc1833              :in std_logic_vector(8 DOWNTO 0);
     Lc1834              :in std_logic_vector(8 DOWNTO 0);
     Lc1835              :in std_logic_vector(8 DOWNTO 0);
     Lc1836              :in std_logic_vector(8 DOWNTO 0);
     Lc1837              :in std_logic_vector(8 DOWNTO 0);
     Lc1838              :in std_logic_vector(8 DOWNTO 0);
     Lc1839              :in std_logic_vector(8 DOWNTO 0);
     Lc1840              :in std_logic_vector(8 DOWNTO 0);
     Lc1841              :in std_logic_vector(8 DOWNTO 0);
     Lc1842              :in std_logic_vector(8 DOWNTO 0);
     Lc1843              :in std_logic_vector(8 DOWNTO 0);
     Lc1844              :in std_logic_vector(8 DOWNTO 0);
     Lc1845              :in std_logic_vector(8 DOWNTO 0);
     Lc1846              :in std_logic_vector(8 DOWNTO 0);
     Lc1847              :in std_logic_vector(8 DOWNTO 0);
     Lc1848              :in std_logic_vector(8 DOWNTO 0);
     Lc1849              :in std_logic_vector(8 DOWNTO 0);
     Lc1850              :in std_logic_vector(8 DOWNTO 0);
     Lc1851              :in std_logic_vector(8 DOWNTO 0);
     Lc1852              :in std_logic_vector(8 DOWNTO 0);
     Lc1853              :in std_logic_vector(8 DOWNTO 0);
     Lc1854              :in std_logic_vector(8 DOWNTO 0);
     Lc1855              :in std_logic_vector(8 DOWNTO 0);
     Lc1856              :in std_logic_vector(8 DOWNTO 0);
     Lc1857              :in std_logic_vector(8 DOWNTO 0);
     Lc1858              :in std_logic_vector(8 DOWNTO 0);
     Lc1859              :in std_logic_vector(8 DOWNTO 0);
     Lc1860              :in std_logic_vector(8 DOWNTO 0);
     Lc1861              :in std_logic_vector(8 DOWNTO 0);
     Lc1862              :in std_logic_vector(8 DOWNTO 0);
     Lc1863              :in std_logic_vector(8 DOWNTO 0);
     Lc1864              :in std_logic_vector(8 DOWNTO 0);
     Lc1865              :in std_logic_vector(8 DOWNTO 0);
     Lc1866              :in std_logic_vector(8 DOWNTO 0);
     Lc1867              :in std_logic_vector(8 DOWNTO 0);
     Lc1868              :in std_logic_vector(8 DOWNTO 0);
     Lc1869              :in std_logic_vector(8 DOWNTO 0);
     Lc1870              :in std_logic_vector(8 DOWNTO 0);
     Lc1871              :in std_logic_vector(8 DOWNTO 0);
     Lc1872              :in std_logic_vector(8 DOWNTO 0);
     Lc1873              :in std_logic_vector(8 DOWNTO 0);
     Lc1874              :in std_logic_vector(8 DOWNTO 0);
     Lc1875              :in std_logic_vector(8 DOWNTO 0);
     Lc1876              :in std_logic_vector(8 DOWNTO 0);
     Lc1877              :in std_logic_vector(8 DOWNTO 0);
     Lc1878              :in std_logic_vector(8 DOWNTO 0);
     Lc1879              :in std_logic_vector(8 DOWNTO 0);
     Lc1880              :in std_logic_vector(8 DOWNTO 0);
     Lc1881              :in std_logic_vector(8 DOWNTO 0);
     Lc1882              :in std_logic_vector(8 DOWNTO 0);
     Lc1883              :in std_logic_vector(8 DOWNTO 0);
     Lc1884              :in std_logic_vector(8 DOWNTO 0);
     Lc1885              :in std_logic_vector(8 DOWNTO 0);
     Lc1886              :in std_logic_vector(8 DOWNTO 0);
     Lc1887              :in std_logic_vector(8 DOWNTO 0);
     Lc1888              :in std_logic_vector(8 DOWNTO 0);
     Lc1889              :in std_logic_vector(8 DOWNTO 0);
     Lc1890              :in std_logic_vector(8 DOWNTO 0);
     Lc1891              :in std_logic_vector(8 DOWNTO 0);
     Lc1892              :in std_logic_vector(8 DOWNTO 0);
     Lc1893              :in std_logic_vector(8 DOWNTO 0);
     Lc1894              :in std_logic_vector(8 DOWNTO 0);
     Lc1895              :in std_logic_vector(8 DOWNTO 0);
     Lc1896              :in std_logic_vector(8 DOWNTO 0);
     Lc1897              :in std_logic_vector(8 DOWNTO 0);
     Lc1898              :in std_logic_vector(8 DOWNTO 0);
     Lc1899              :in std_logic_vector(8 DOWNTO 0);
     Lc1900              :in std_logic_vector(8 DOWNTO 0);
     Lc1901              :in std_logic_vector(8 DOWNTO 0);
     Lc1902              :in std_logic_vector(8 DOWNTO 0);
     Lc1903              :in std_logic_vector(8 DOWNTO 0);
     Lc1904              :in std_logic_vector(8 DOWNTO 0);
     Lc1905              :in std_logic_vector(8 DOWNTO 0);
     Lc1906              :in std_logic_vector(8 DOWNTO 0);
     Lc1907              :in std_logic_vector(8 DOWNTO 0);
     Lc1908              :in std_logic_vector(8 DOWNTO 0);
     Lc1909              :in std_logic_vector(8 DOWNTO 0);
     Lc1910              :in std_logic_vector(8 DOWNTO 0);
     Lc1911              :in std_logic_vector(8 DOWNTO 0);
     Lc1912              :in std_logic_vector(8 DOWNTO 0);
     Lc1913              :in std_logic_vector(8 DOWNTO 0);
     Lc1914              :in std_logic_vector(8 DOWNTO 0);
     Lc1915              :in std_logic_vector(8 DOWNTO 0);
     Lc1916              :in std_logic_vector(8 DOWNTO 0);
     Lc1917              :in std_logic_vector(8 DOWNTO 0);
     Lc1918              :in std_logic_vector(8 DOWNTO 0);
     Lc1919              :in std_logic_vector(8 DOWNTO 0);
     Lc1920              :in std_logic_vector(8 DOWNTO 0);
     Lc1921              :in std_logic_vector(8 DOWNTO 0);
     Lc1922              :in std_logic_vector(8 DOWNTO 0);
     Lc1923              :in std_logic_vector(8 DOWNTO 0);
     Lc1924              :in std_logic_vector(8 DOWNTO 0);
     Lc1925              :in std_logic_vector(8 DOWNTO 0);
     Lc1926              :in std_logic_vector(8 DOWNTO 0);
     Lc1927              :in std_logic_vector(8 DOWNTO 0);
     Lc1928              :in std_logic_vector(8 DOWNTO 0);
     Lc1929              :in std_logic_vector(8 DOWNTO 0);
     Lc1930              :in std_logic_vector(8 DOWNTO 0);
     Lc1931              :in std_logic_vector(8 DOWNTO 0);
     Lc1932              :in std_logic_vector(8 DOWNTO 0);
     Lc1933              :in std_logic_vector(8 DOWNTO 0);
     Lc1934              :in std_logic_vector(8 DOWNTO 0);
     Lc1935              :in std_logic_vector(8 DOWNTO 0);
     Lc1936              :in std_logic_vector(8 DOWNTO 0);
     Lc1937              :in std_logic_vector(8 DOWNTO 0);
     Lc1938              :in std_logic_vector(8 DOWNTO 0);
     Lc1939              :in std_logic_vector(8 DOWNTO 0);
     Lc1940              :in std_logic_vector(8 DOWNTO 0);
     Lc1941              :in std_logic_vector(8 DOWNTO 0);
     Lc1942              :in std_logic_vector(8 DOWNTO 0);
     Lc1943              :in std_logic_vector(8 DOWNTO 0);
     Lc1944              :in std_logic_vector(8 DOWNTO 0);
     Lc1945              :in std_logic_vector(8 DOWNTO 0);
     Lc1946              :in std_logic_vector(8 DOWNTO 0);
     Lc1947              :in std_logic_vector(8 DOWNTO 0);
     Lc1948              :in std_logic_vector(8 DOWNTO 0);
     Lc1949              :in std_logic_vector(8 DOWNTO 0);
     Lc1950              :in std_logic_vector(8 DOWNTO 0);
     Lc1951              :in std_logic_vector(8 DOWNTO 0);
     Lc1952              :in std_logic_vector(8 DOWNTO 0);
     Lc1953              :in std_logic_vector(8 DOWNTO 0);
     Lc1954              :in std_logic_vector(8 DOWNTO 0);
     Lc1955              :in std_logic_vector(8 DOWNTO 0);
     Lc1956              :in std_logic_vector(8 DOWNTO 0);
     Lc1957              :in std_logic_vector(8 DOWNTO 0);
     Lc1958              :in std_logic_vector(8 DOWNTO 0);
     Lc1959              :in std_logic_vector(8 DOWNTO 0);
     Lc1960              :in std_logic_vector(8 DOWNTO 0);
     Lc1961              :in std_logic_vector(8 DOWNTO 0);
     Lc1962              :in std_logic_vector(8 DOWNTO 0);
     Lc1963              :in std_logic_vector(8 DOWNTO 0);
     Lc1964              :in std_logic_vector(8 DOWNTO 0);
     Lc1965              :in std_logic_vector(8 DOWNTO 0);
     Lc1966              :in std_logic_vector(8 DOWNTO 0);
     Lc1967              :in std_logic_vector(8 DOWNTO 0);
     Lc1968              :in std_logic_vector(8 DOWNTO 0);
     Lc1969              :in std_logic_vector(8 DOWNTO 0);
     Lc1970              :in std_logic_vector(8 DOWNTO 0);
     Lc1971              :in std_logic_vector(8 DOWNTO 0);
     Lc1972              :in std_logic_vector(8 DOWNTO 0);
     Lc1973              :in std_logic_vector(8 DOWNTO 0);
     Lc1974              :in std_logic_vector(8 DOWNTO 0);
     Lc1975              :in std_logic_vector(8 DOWNTO 0);
     Lc1976              :in std_logic_vector(8 DOWNTO 0);
     Lc1977              :in std_logic_vector(8 DOWNTO 0);
     Lc1978              :in std_logic_vector(8 DOWNTO 0);
     Lc1979              :in std_logic_vector(8 DOWNTO 0);
     Lc1980              :in std_logic_vector(8 DOWNTO 0);
     Lc1981              :in std_logic_vector(8 DOWNTO 0);
     Lc1982              :in std_logic_vector(8 DOWNTO 0);
     Lc1983              :in std_logic_vector(8 DOWNTO 0);
     Lc1984              :in std_logic_vector(8 DOWNTO 0);
     Lc1985              :in std_logic_vector(8 DOWNTO 0);
     Lc1986              :in std_logic_vector(8 DOWNTO 0);
     Lc1987              :in std_logic_vector(8 DOWNTO 0);
     Lc1988              :in std_logic_vector(8 DOWNTO 0);
     Lc1989              :in std_logic_vector(8 DOWNTO 0);
     Lc1990              :in std_logic_vector(8 DOWNTO 0);
     Lc1991              :in std_logic_vector(8 DOWNTO 0);
     Lc1992              :in std_logic_vector(8 DOWNTO 0);
     Lc1993              :in std_logic_vector(8 DOWNTO 0);
     Lc1994              :in std_logic_vector(8 DOWNTO 0);
     Lc1995              :in std_logic_vector(8 DOWNTO 0);
     Lc1996              :in std_logic_vector(8 DOWNTO 0);
     Lc1997              :in std_logic_vector(8 DOWNTO 0);
     Lc1998              :in std_logic_vector(8 DOWNTO 0);
     Lc1999              :in std_logic_vector(8 DOWNTO 0);
     Lc2000              :in std_logic_vector(8 DOWNTO 0);
     Lc2001              :in std_logic_vector(8 DOWNTO 0);
     Lc2002              :in std_logic_vector(8 DOWNTO 0);
     Lc2003              :in std_logic_vector(8 DOWNTO 0);
     Lc2004              :in std_logic_vector(8 DOWNTO 0);
     Lc2005              :in std_logic_vector(8 DOWNTO 0);
     Lc2006              :in std_logic_vector(8 DOWNTO 0);
     Lc2007              :in std_logic_vector(8 DOWNTO 0);
     Lc2008              :in std_logic_vector(8 DOWNTO 0);
     Lc2009              :in std_logic_vector(8 DOWNTO 0);
     Lc2010              :in std_logic_vector(8 DOWNTO 0);
     Lc2011              :in std_logic_vector(8 DOWNTO 0);
     Lc2012              :in std_logic_vector(8 DOWNTO 0);
     Lc2013              :in std_logic_vector(8 DOWNTO 0);
     Lc2014              :in std_logic_vector(8 DOWNTO 0);
     Lc2015              :in std_logic_vector(8 DOWNTO 0);
     Lc2016              :in std_logic_vector(8 DOWNTO 0);
     Lc2017              :in std_logic_vector(8 DOWNTO 0);
     Lc2018              :in std_logic_vector(8 DOWNTO 0);
     Lc2019              :in std_logic_vector(8 DOWNTO 0);
     Lc2020              :in std_logic_vector(8 DOWNTO 0);
     Lc2021              :in std_logic_vector(8 DOWNTO 0);
     Lc2022              :in std_logic_vector(8 DOWNTO 0);
     Lc2023              :in std_logic_vector(8 DOWNTO 0);
     Lc2024              :in std_logic_vector(8 DOWNTO 0);
     Lc2025              :in std_logic_vector(8 DOWNTO 0);
     Lc2026              :in std_logic_vector(8 DOWNTO 0);
     Lc2027              :in std_logic_vector(8 DOWNTO 0);
     Lc2028              :in std_logic_vector(8 DOWNTO 0);
     Lc2029              :in std_logic_vector(8 DOWNTO 0);
     Lc2030              :in std_logic_vector(8 DOWNTO 0);
     Lc2031              :in std_logic_vector(8 DOWNTO 0);
     Lc2032              :in std_logic_vector(8 DOWNTO 0);
     Lc2033              :in std_logic_vector(8 DOWNTO 0);
     Lc2034              :in std_logic_vector(8 DOWNTO 0);
     Lc2035              :in std_logic_vector(8 DOWNTO 0);
     Lc2036              :in std_logic_vector(8 DOWNTO 0);
     Lc2037              :in std_logic_vector(8 DOWNTO 0);
     Lc2038              :in std_logic_vector(8 DOWNTO 0);
     Lc2039              :in std_logic_vector(8 DOWNTO 0);
     Lc2040              :in std_logic_vector(8 DOWNTO 0);
     Lc2041              :in std_logic_vector(8 DOWNTO 0);
     Lc2042              :in std_logic_vector(8 DOWNTO 0);
     Lc2043              :in std_logic_vector(8 DOWNTO 0);
     Lc2044              :in std_logic_vector(8 DOWNTO 0);
     Lc2045              :in std_logic_vector(8 DOWNTO 0);
     Lc2046              :in std_logic_vector(8 DOWNTO 0);
     Lc2047              :in std_logic_vector(8 DOWNTO 0);
     Lc2048              :in std_logic_vector(8 DOWNTO 0);
     Lc2049              :in std_logic_vector(8 DOWNTO 0);
     Lc2050              :in std_logic_vector(8 DOWNTO 0);
     Lc2051              :in std_logic_vector(8 DOWNTO 0);
     Lc2052              :in std_logic_vector(8 DOWNTO 0);
     Lc2053              :in std_logic_vector(8 DOWNTO 0);
     Lc2054              :in std_logic_vector(8 DOWNTO 0);
     Lc2055              :in std_logic_vector(8 DOWNTO 0);
     Lc2056              :in std_logic_vector(8 DOWNTO 0);
     Lc2057              :in std_logic_vector(8 DOWNTO 0);
     Lc2058              :in std_logic_vector(8 DOWNTO 0);
     Lc2059              :in std_logic_vector(8 DOWNTO 0);
     Lc2060              :in std_logic_vector(8 DOWNTO 0);
     Lc2061              :in std_logic_vector(8 DOWNTO 0);
     Lc2062              :in std_logic_vector(8 DOWNTO 0);
     Lc2063              :in std_logic_vector(8 DOWNTO 0);
     Lc2064              :in std_logic_vector(8 DOWNTO 0);
     Lc2065              :in std_logic_vector(8 DOWNTO 0);
     Lc2066              :in std_logic_vector(8 DOWNTO 0);
     Lc2067              :in std_logic_vector(8 DOWNTO 0);
     Lc2068              :in std_logic_vector(8 DOWNTO 0);
     Lc2069              :in std_logic_vector(8 DOWNTO 0);
     Lc2070              :in std_logic_vector(8 DOWNTO 0);
     Lc2071              :in std_logic_vector(8 DOWNTO 0);
     Lc2072              :in std_logic_vector(8 DOWNTO 0);
     Lc2073              :in std_logic_vector(8 DOWNTO 0);
     Lc2074              :in std_logic_vector(8 DOWNTO 0);
     Lc2075              :in std_logic_vector(8 DOWNTO 0);
     Lc2076              :in std_logic_vector(8 DOWNTO 0);
     Lc2077              :in std_logic_vector(8 DOWNTO 0);
     Lc2078              :in std_logic_vector(8 DOWNTO 0);
     Lc2079              :in std_logic_vector(8 DOWNTO 0);
     Lc2080              :in std_logic_vector(8 DOWNTO 0);
     Lc2081              :in std_logic_vector(8 DOWNTO 0);
     Lc2082              :in std_logic_vector(8 DOWNTO 0);
     Lc2083              :in std_logic_vector(8 DOWNTO 0);
     Lc2084              :in std_logic_vector(8 DOWNTO 0);
     Lc2085              :in std_logic_vector(8 DOWNTO 0);
     Lc2086              :in std_logic_vector(8 DOWNTO 0);
     Lc2087              :in std_logic_vector(8 DOWNTO 0);
     Lc2088              :in std_logic_vector(8 DOWNTO 0);
     Lc2089              :in std_logic_vector(8 DOWNTO 0);
     Lc2090              :in std_logic_vector(8 DOWNTO 0);
     Lc2091              :in std_logic_vector(8 DOWNTO 0);
     Lc2092              :in std_logic_vector(8 DOWNTO 0);
     Lc2093              :in std_logic_vector(8 DOWNTO 0);
     Lc2094              :in std_logic_vector(8 DOWNTO 0);
     Lc2095              :in std_logic_vector(8 DOWNTO 0);
     Lc2096              :in std_logic_vector(8 DOWNTO 0);
     Lc2097              :in std_logic_vector(8 DOWNTO 0);
     Lc2098              :in std_logic_vector(8 DOWNTO 0);
     Lc2099              :in std_logic_vector(8 DOWNTO 0);
     Lc2100              :in std_logic_vector(8 DOWNTO 0);
     Lc2101              :in std_logic_vector(8 DOWNTO 0);
     Lc2102              :in std_logic_vector(8 DOWNTO 0);
     Lc2103              :in std_logic_vector(8 DOWNTO 0);
     Lc2104              :in std_logic_vector(8 DOWNTO 0);
     Lc2105              :in std_logic_vector(8 DOWNTO 0);
     Lc2106              :in std_logic_vector(8 DOWNTO 0);
     Lc2107              :in std_logic_vector(8 DOWNTO 0);
     Lc2108              :in std_logic_vector(8 DOWNTO 0);
     Lc2109              :in std_logic_vector(8 DOWNTO 0);
     Lc2110              :in std_logic_vector(8 DOWNTO 0);
     Lc2111              :in std_logic_vector(8 DOWNTO 0);
     Lc2112              :in std_logic_vector(8 DOWNTO 0);
     Lc2113              :in std_logic_vector(8 DOWNTO 0);
     Lc2114              :in std_logic_vector(8 DOWNTO 0);
     Lc2115              :in std_logic_vector(8 DOWNTO 0);
     Lc2116              :in std_logic_vector(8 DOWNTO 0);
     Lc2117              :in std_logic_vector(8 DOWNTO 0);
     Lc2118              :in std_logic_vector(8 DOWNTO 0);
     Lc2119              :in std_logic_vector(8 DOWNTO 0);
     Lc2120              :in std_logic_vector(8 DOWNTO 0);
     Lc2121              :in std_logic_vector(8 DOWNTO 0);
     Lc2122              :in std_logic_vector(8 DOWNTO 0);
     Lc2123              :in std_logic_vector(8 DOWNTO 0);
     Lc2124              :in std_logic_vector(8 DOWNTO 0);
     Lc2125              :in std_logic_vector(8 DOWNTO 0);
     Lc2126              :in std_logic_vector(8 DOWNTO 0);
     Lc2127              :in std_logic_vector(8 DOWNTO 0);
     Lc2128              :in std_logic_vector(8 DOWNTO 0);
     Lc2129              :in std_logic_vector(8 DOWNTO 0);
     Lc2130              :in std_logic_vector(8 DOWNTO 0);
     Lc2131              :in std_logic_vector(8 DOWNTO 0);
     Lc2132              :in std_logic_vector(8 DOWNTO 0);
     Lc2133              :in std_logic_vector(8 DOWNTO 0);
     Lc2134              :in std_logic_vector(8 DOWNTO 0);
     Lc2135              :in std_logic_vector(8 DOWNTO 0);
     Lc2136              :in std_logic_vector(8 DOWNTO 0);
     Lc2137              :in std_logic_vector(8 DOWNTO 0);
     Lc2138              :in std_logic_vector(8 DOWNTO 0);
     Lc2139              :in std_logic_vector(8 DOWNTO 0);
     Lc2140              :in std_logic_vector(8 DOWNTO 0);
     Lc2141              :in std_logic_vector(8 DOWNTO 0);
     Lc2142              :in std_logic_vector(8 DOWNTO 0);
     Lc2143              :in std_logic_vector(8 DOWNTO 0);
     Lc2144              :in std_logic_vector(8 DOWNTO 0);
     Lc2145              :in std_logic_vector(8 DOWNTO 0);
     Lc2146              :in std_logic_vector(8 DOWNTO 0);
     Lc2147              :in std_logic_vector(8 DOWNTO 0);
     Lc2148              :in std_logic_vector(8 DOWNTO 0);
     Lc2149              :in std_logic_vector(8 DOWNTO 0);
     Lc2150              :in std_logic_vector(8 DOWNTO 0);
     Lc2151              :in std_logic_vector(8 DOWNTO 0);
     Lc2152              :in std_logic_vector(8 DOWNTO 0);
     Lc2153              :in std_logic_vector(8 DOWNTO 0);
     Lc2154              :in std_logic_vector(8 DOWNTO 0);
     Lc2155              :in std_logic_vector(8 DOWNTO 0);
     Lc2156              :in std_logic_vector(8 DOWNTO 0);
     Lc2157              :in std_logic_vector(8 DOWNTO 0);
     Lc2158              :in std_logic_vector(8 DOWNTO 0);
     Lc2159              :in std_logic_vector(8 DOWNTO 0);
     Lc2160              :in std_logic_vector(8 DOWNTO 0);
     Lc2161              :in std_logic_vector(8 DOWNTO 0);
     Lc2162              :in std_logic_vector(8 DOWNTO 0);
     Lc2163              :in std_logic_vector(8 DOWNTO 0);
     Lc2164              :in std_logic_vector(8 DOWNTO 0);
     Lc2165              :in std_logic_vector(8 DOWNTO 0);
     Lc2166              :in std_logic_vector(8 DOWNTO 0);
     Lc2167              :in std_logic_vector(8 DOWNTO 0);
     Lc2168              :in std_logic_vector(8 DOWNTO 0);
     Lc2169              :in std_logic_vector(8 DOWNTO 0);
     Lc2170              :in std_logic_vector(8 DOWNTO 0);
     Lc2171              :in std_logic_vector(8 DOWNTO 0);
     Lc2172              :in std_logic_vector(8 DOWNTO 0);
     Lc2173              :in std_logic_vector(8 DOWNTO 0);
     Lc2174              :in std_logic_vector(8 DOWNTO 0);
     Lc2175              :in std_logic_vector(8 DOWNTO 0);
     Lc2176              :in std_logic_vector(8 DOWNTO 0);
     Lc2177              :in std_logic_vector(8 DOWNTO 0);
     Lc2178              :in std_logic_vector(8 DOWNTO 0);
     Lc2179              :in std_logic_vector(8 DOWNTO 0);
     Lc2180              :in std_logic_vector(8 DOWNTO 0);
     Lc2181              :in std_logic_vector(8 DOWNTO 0);
     Lc2182              :in std_logic_vector(8 DOWNTO 0);
     Lc2183              :in std_logic_vector(8 DOWNTO 0);
     Lc2184              :in std_logic_vector(8 DOWNTO 0);
     Lc2185              :in std_logic_vector(8 DOWNTO 0);
     Lc2186              :in std_logic_vector(8 DOWNTO 0);
     Lc2187              :in std_logic_vector(8 DOWNTO 0);
     Lc2188              :in std_logic_vector(8 DOWNTO 0);
     Lc2189              :in std_logic_vector(8 DOWNTO 0);
     Lc2190              :in std_logic_vector(8 DOWNTO 0);
     Lc2191              :in std_logic_vector(8 DOWNTO 0);
     Lc2192              :in std_logic_vector(8 DOWNTO 0);
     Lc2193              :in std_logic_vector(8 DOWNTO 0);
     Lc2194              :in std_logic_vector(8 DOWNTO 0);
     Lc2195              :in std_logic_vector(8 DOWNTO 0);
     Lc2196              :in std_logic_vector(8 DOWNTO 0);
     Lc2197              :in std_logic_vector(8 DOWNTO 0);
     Lc2198              :in std_logic_vector(8 DOWNTO 0);
     Lc2199              :in std_logic_vector(8 DOWNTO 0);
     Lc2200              :in std_logic_vector(8 DOWNTO 0);
     Lc2201              :in std_logic_vector(8 DOWNTO 0);
     Lc2202              :in std_logic_vector(8 DOWNTO 0);
     Lc2203              :in std_logic_vector(8 DOWNTO 0);
     Lc2204              :in std_logic_vector(8 DOWNTO 0);
     Lc2205              :in std_logic_vector(8 DOWNTO 0);
     Lc2206              :in std_logic_vector(8 DOWNTO 0);
     Lc2207              :in std_logic_vector(8 DOWNTO 0);
     Lc2208              :in std_logic_vector(8 DOWNTO 0);
     Lc2209              :in std_logic_vector(8 DOWNTO 0);
     Lc2210              :in std_logic_vector(8 DOWNTO 0);
     Lc2211              :in std_logic_vector(8 DOWNTO 0);
     Lc2212              :in std_logic_vector(8 DOWNTO 0);
     Lc2213              :in std_logic_vector(8 DOWNTO 0);
     Lc2214              :in std_logic_vector(8 DOWNTO 0);
     Lc2215              :in std_logic_vector(8 DOWNTO 0);
     Lc2216              :in std_logic_vector(8 DOWNTO 0);
     Lc2217              :in std_logic_vector(8 DOWNTO 0);
     Lc2218              :in std_logic_vector(8 DOWNTO 0);
     Lc2219              :in std_logic_vector(8 DOWNTO 0);
     Lc2220              :in std_logic_vector(8 DOWNTO 0);
     Lc2221              :in std_logic_vector(8 DOWNTO 0);
     Lc2222              :in std_logic_vector(8 DOWNTO 0);
     Lc2223              :in std_logic_vector(8 DOWNTO 0);
     Lc2224              :in std_logic_vector(8 DOWNTO 0);
     Lc2225              :in std_logic_vector(8 DOWNTO 0);
     Lc2226              :in std_logic_vector(8 DOWNTO 0);
     Lc2227              :in std_logic_vector(8 DOWNTO 0);
     Lc2228              :in std_logic_vector(8 DOWNTO 0);
     Lc2229              :in std_logic_vector(8 DOWNTO 0);
     Lc2230              :in std_logic_vector(8 DOWNTO 0);
     Lc2231              :in std_logic_vector(8 DOWNTO 0);
     Lc2232              :in std_logic_vector(8 DOWNTO 0);
     Lc2233              :in std_logic_vector(8 DOWNTO 0);
     Lc2234              :in std_logic_vector(8 DOWNTO 0);
     Lc2235              :in std_logic_vector(8 DOWNTO 0);
     Lc2236              :in std_logic_vector(8 DOWNTO 0);
     Lc2237              :in std_logic_vector(8 DOWNTO 0);
     Lc2238              :in std_logic_vector(8 DOWNTO 0);
     Lc2239              :in std_logic_vector(8 DOWNTO 0);
     Lc2240              :in std_logic_vector(8 DOWNTO 0);
     Lc2241              :in std_logic_vector(8 DOWNTO 0);
     Lc2242              :in std_logic_vector(8 DOWNTO 0);
     Lc2243              :in std_logic_vector(8 DOWNTO 0);
     Lc2244              :in std_logic_vector(8 DOWNTO 0);
     Lc2245              :in std_logic_vector(8 DOWNTO 0);
     Lc2246              :in std_logic_vector(8 DOWNTO 0);
     Lc2247              :in std_logic_vector(8 DOWNTO 0);
     Lc2248              :in std_logic_vector(8 DOWNTO 0);
     Lc2249              :in std_logic_vector(8 DOWNTO 0);
     Lc2250              :in std_logic_vector(8 DOWNTO 0);
     Lc2251              :in std_logic_vector(8 DOWNTO 0);
     Lc2252              :in std_logic_vector(8 DOWNTO 0);
     Lc2253              :in std_logic_vector(8 DOWNTO 0);
     Lc2254              :in std_logic_vector(8 DOWNTO 0);
     Lc2255              :in std_logic_vector(8 DOWNTO 0);
     Lc2256              :in std_logic_vector(8 DOWNTO 0);
     Lc2257              :in std_logic_vector(8 DOWNTO 0);
     Lc2258              :in std_logic_vector(8 DOWNTO 0);
     Lc2259              :in std_logic_vector(8 DOWNTO 0);
     Lc2260              :in std_logic_vector(8 DOWNTO 0);
     Lc2261              :in std_logic_vector(8 DOWNTO 0);
     Lc2262              :in std_logic_vector(8 DOWNTO 0);
     Lc2263              :in std_logic_vector(8 DOWNTO 0);
     Lc2264              :in std_logic_vector(8 DOWNTO 0);
     Lc2265              :in std_logic_vector(8 DOWNTO 0);
     Lc2266              :in std_logic_vector(8 DOWNTO 0);
     Lc2267              :in std_logic_vector(8 DOWNTO 0);
     Lc2268              :in std_logic_vector(8 DOWNTO 0);
     Lc2269              :in std_logic_vector(8 DOWNTO 0);
     Lc2270              :in std_logic_vector(8 DOWNTO 0);
     Lc2271              :in std_logic_vector(8 DOWNTO 0);
     Lc2272              :in std_logic_vector(8 DOWNTO 0);
     Lc2273              :in std_logic_vector(8 DOWNTO 0);
     Lc2274              :in std_logic_vector(8 DOWNTO 0);
     Lc2275              :in std_logic_vector(8 DOWNTO 0);
     Lc2276              :in std_logic_vector(8 DOWNTO 0);
     Lc2277              :in std_logic_vector(8 DOWNTO 0);
     Lc2278              :in std_logic_vector(8 DOWNTO 0);
     Lc2279              :in std_logic_vector(8 DOWNTO 0);
     Lc2280              :in std_logic_vector(8 DOWNTO 0);
     Lc2281              :in std_logic_vector(8 DOWNTO 0);
     Lc2282              :in std_logic_vector(8 DOWNTO 0);
     Lc2283              :in std_logic_vector(8 DOWNTO 0);
     Lc2284              :in std_logic_vector(8 DOWNTO 0);
     Lc2285              :in std_logic_vector(8 DOWNTO 0);
     Lc2286              :in std_logic_vector(8 DOWNTO 0);
     Lc2287              :in std_logic_vector(8 DOWNTO 0);
     Lc2288              :in std_logic_vector(8 DOWNTO 0);
     Lc2289              :in std_logic_vector(8 DOWNTO 0);
     Lc2290              :in std_logic_vector(8 DOWNTO 0);
     Lc2291              :in std_logic_vector(8 DOWNTO 0);
     Lc2292              :in std_logic_vector(8 DOWNTO 0);
     Lc2293              :in std_logic_vector(8 DOWNTO 0);
     Lc2294              :in std_logic_vector(8 DOWNTO 0);
     Lc2295              :in std_logic_vector(8 DOWNTO 0);
     Lc2296              :in std_logic_vector(8 DOWNTO 0);
     Lc2297              :in std_logic_vector(8 DOWNTO 0);
     Lc2298              :in std_logic_vector(8 DOWNTO 0);
     Lc2299              :in std_logic_vector(8 DOWNTO 0);
     Lc2300              :in std_logic_vector(8 DOWNTO 0);
     Lc2301              :in std_logic_vector(8 DOWNTO 0);
     Lc2302              :in std_logic_vector(8 DOWNTO 0);
     Lc2303              :in std_logic_vector(8 DOWNTO 0);
     Lc2304              :in std_logic_vector(8 DOWNTO 0);
     out1            :out std_logic;
     out2            :out std_logic;
     out3            :out std_logic;
     out4            :out std_logic;
     out5            :out std_logic;
     out6            :out std_logic;
     out7            :out std_logic;
     out8            :out std_logic;
     out9            :out std_logic;
     out10            :out std_logic;
     out11            :out std_logic;
     out12            :out std_logic;
     out13            :out std_logic;
     out14            :out std_logic;
     out15            :out std_logic;
     out16            :out std_logic;
     out17            :out std_logic;
     out18            :out std_logic;
     out19            :out std_logic;
     out20            :out std_logic;
     out21            :out std_logic;
     out22            :out std_logic;
     out23            :out std_logic;
     out24            :out std_logic;
     out25            :out std_logic;
     out26            :out std_logic;
     out27            :out std_logic;
     out28            :out std_logic;
     out29            :out std_logic;
     out30            :out std_logic;
     out31            :out std_logic;
     out32            :out std_logic;
     out33            :out std_logic;
     out34            :out std_logic;
     out35            :out std_logic;
     out36            :out std_logic;
     out37            :out std_logic;
     out38            :out std_logic;
     out39            :out std_logic;
     out40            :out std_logic;
     out41            :out std_logic;
     out42            :out std_logic;
     out43            :out std_logic;
     out44            :out std_logic;
     out45            :out std_logic;
     out46            :out std_logic;
     out47            :out std_logic;
     out48            :out std_logic;
     out49            :out std_logic;
     out50            :out std_logic;
     out51            :out std_logic;
     out52            :out std_logic;
     out53            :out std_logic;
     out54            :out std_logic;
     out55            :out std_logic;
     out56            :out std_logic;
     out57            :out std_logic;
     out58            :out std_logic;
     out59            :out std_logic;
     out60            :out std_logic;
     out61            :out std_logic;
     out62            :out std_logic;
     out63            :out std_logic;
     out64            :out std_logic;
     out65            :out std_logic;
     out66            :out std_logic;
     out67            :out std_logic;
     out68            :out std_logic;
     out69            :out std_logic;
     out70            :out std_logic;
     out71            :out std_logic;
     out72            :out std_logic;
     out73            :out std_logic;
     out74            :out std_logic;
     out75            :out std_logic;
     out76            :out std_logic;
     out77            :out std_logic;
     out78            :out std_logic;
     out79            :out std_logic;
     out80            :out std_logic;
     out81            :out std_logic;
     out82            :out std_logic;
     out83            :out std_logic;
     out84            :out std_logic;
     out85            :out std_logic;
     out86            :out std_logic;
     out87            :out std_logic;
     out88            :out std_logic;
     out89            :out std_logic;
     out90            :out std_logic;
     out91            :out std_logic;
     out92            :out std_logic;
     out93            :out std_logic;
     out94            :out std_logic;
     out95            :out std_logic;
     out96            :out std_logic;
     out97            :out std_logic;
     out98            :out std_logic;
     out99            :out std_logic;
     out100            :out std_logic;
     out101            :out std_logic;
     out102            :out std_logic;
     out103            :out std_logic;
     out104            :out std_logic;
     out105            :out std_logic;
     out106            :out std_logic;
     out107            :out std_logic;
     out108            :out std_logic;
     out109            :out std_logic;
     out110            :out std_logic;
     out111            :out std_logic;
     out112            :out std_logic;
     out113            :out std_logic;
     out114            :out std_logic;
     out115            :out std_logic;
     out116            :out std_logic;
     out117            :out std_logic;
     out118            :out std_logic;
     out119            :out std_logic;
     out120            :out std_logic;
     out121            :out std_logic;
     out122            :out std_logic;
     out123            :out std_logic;
     out124            :out std_logic;
     out125            :out std_logic;
     out126            :out std_logic;
     out127            :out std_logic;
     out128            :out std_logic;
     out129            :out std_logic;
     out130            :out std_logic;
     out131            :out std_logic;
     out132            :out std_logic;
     out133            :out std_logic;
     out134            :out std_logic;
     out135            :out std_logic;
     out136            :out std_logic;
     out137            :out std_logic;
     out138            :out std_logic;
     out139            :out std_logic;
     out140            :out std_logic;
     out141            :out std_logic;
     out142            :out std_logic;
     out143            :out std_logic;
     out144            :out std_logic;
     out145            :out std_logic;
     out146            :out std_logic;
     out147            :out std_logic;
     out148            :out std_logic;
     out149            :out std_logic;
     out150            :out std_logic;
     out151            :out std_logic;
     out152            :out std_logic;
     out153            :out std_logic;
     out154            :out std_logic;
     out155            :out std_logic;
     out156            :out std_logic;
     out157            :out std_logic;
     out158            :out std_logic;
     out159            :out std_logic;
     out160            :out std_logic;
     out161            :out std_logic;
     out162            :out std_logic;
     out163            :out std_logic;
     out164            :out std_logic;
     out165            :out std_logic;
     out166            :out std_logic;
     out167            :out std_logic;
     out168            :out std_logic;
     out169            :out std_logic;
     out170            :out std_logic;
     out171            :out std_logic;
     out172            :out std_logic;
     out173            :out std_logic;
     out174            :out std_logic;
     out175            :out std_logic;
     out176            :out std_logic;
     out177            :out std_logic;
     out178            :out std_logic;
     out179            :out std_logic;
     out180            :out std_logic;
     out181            :out std_logic;
     out182            :out std_logic;
     out183            :out std_logic;
     out184            :out std_logic;
     out185            :out std_logic;
     out186            :out std_logic;
     out187            :out std_logic;
     out188            :out std_logic;
     out189            :out std_logic;
     out190            :out std_logic;
     out191            :out std_logic;
     out192            :out std_logic;
     out193            :out std_logic;
     out194            :out std_logic;
     out195            :out std_logic;
     out196            :out std_logic;
     out197            :out std_logic;
     out198            :out std_logic;
     out199            :out std_logic;
     out200            :out std_logic;
     out201            :out std_logic;
     out202            :out std_logic;
     out203            :out std_logic;
     out204            :out std_logic;
     out205            :out std_logic;
     out206            :out std_logic;
     out207            :out std_logic;
     out208            :out std_logic;
     out209            :out std_logic;
     out210            :out std_logic;
     out211            :out std_logic;
     out212            :out std_logic;
     out213            :out std_logic;
     out214            :out std_logic;
     out215            :out std_logic;
     out216            :out std_logic;
     out217            :out std_logic;
     out218            :out std_logic;
     out219            :out std_logic;
     out220            :out std_logic;
     out221            :out std_logic;
     out222            :out std_logic;
     out223            :out std_logic;
     out224            :out std_logic;
     out225            :out std_logic;
     out226            :out std_logic;
     out227            :out std_logic;
     out228            :out std_logic;
     out229            :out std_logic;
     out230            :out std_logic;
     out231            :out std_logic;
     out232            :out std_logic;
     out233            :out std_logic;
     out234            :out std_logic;
     out235            :out std_logic;
     out236            :out std_logic;
     out237            :out std_logic;
     out238            :out std_logic;
     out239            :out std_logic;
     out240            :out std_logic;
     out241            :out std_logic;
     out242            :out std_logic;
     out243            :out std_logic;
     out244            :out std_logic;
     out245            :out std_logic;
     out246            :out std_logic;
     out247            :out std_logic;
     out248            :out std_logic;
     out249            :out std_logic;
     out250            :out std_logic;
     out251            :out std_logic;
     out252            :out std_logic;
     out253            :out std_logic;
     out254            :out std_logic;
     out255            :out std_logic;
     out256            :out std_logic;
     out257            :out std_logic;
     out258            :out std_logic;
     out259            :out std_logic;
     out260            :out std_logic;
     out261            :out std_logic;
     out262            :out std_logic;
     out263            :out std_logic;
     out264            :out std_logic;
     out265            :out std_logic;
     out266            :out std_logic;
     out267            :out std_logic;
     out268            :out std_logic;
     out269            :out std_logic;
     out270            :out std_logic;
     out271            :out std_logic;
     out272            :out std_logic;
     out273            :out std_logic;
     out274            :out std_logic;
     out275            :out std_logic;
     out276            :out std_logic;
     out277            :out std_logic;
     out278            :out std_logic;
     out279            :out std_logic;
     out280            :out std_logic;
     out281            :out std_logic;
     out282            :out std_logic;
     out283            :out std_logic;
     out284            :out std_logic;
     out285            :out std_logic;
     out286            :out std_logic;
     out287            :out std_logic;
     out288            :out std_logic;
     out289            :out std_logic;
     out290            :out std_logic;
     out291            :out std_logic;
     out292            :out std_logic;
     out293            :out std_logic;
     out294            :out std_logic;
     out295            :out std_logic;
     out296            :out std_logic;
     out297            :out std_logic;
     out298            :out std_logic;
     out299            :out std_logic;
     out300            :out std_logic;
     out301            :out std_logic;
     out302            :out std_logic;
     out303            :out std_logic;
     out304            :out std_logic;
     out305            :out std_logic;
     out306            :out std_logic;
     out307            :out std_logic;
     out308            :out std_logic;
     out309            :out std_logic;
     out310            :out std_logic;
     out311            :out std_logic;
     out312            :out std_logic;
     out313            :out std_logic;
     out314            :out std_logic;
     out315            :out std_logic;
     out316            :out std_logic;
     out317            :out std_logic;
     out318            :out std_logic;
     out319            :out std_logic;
     out320            :out std_logic;
     out321            :out std_logic;
     out322            :out std_logic;
     out323            :out std_logic;
     out324            :out std_logic;
     out325            :out std_logic;
     out326            :out std_logic;
     out327            :out std_logic;
     out328            :out std_logic;
     out329            :out std_logic;
     out330            :out std_logic;
     out331            :out std_logic;
     out332            :out std_logic;
     out333            :out std_logic;
     out334            :out std_logic;
     out335            :out std_logic;
     out336            :out std_logic;
     out337            :out std_logic;
     out338            :out std_logic;
     out339            :out std_logic;
     out340            :out std_logic;
     out341            :out std_logic;
     out342            :out std_logic;
     out343            :out std_logic;
     out344            :out std_logic;
     out345            :out std_logic;
     out346            :out std_logic;
     out347            :out std_logic;
     out348            :out std_logic;
     out349            :out std_logic;
     out350            :out std_logic;
     out351            :out std_logic;
     out352            :out std_logic;
     out353            :out std_logic;
     out354            :out std_logic;
     out355            :out std_logic;
     out356            :out std_logic;
     out357            :out std_logic;
     out358            :out std_logic;
     out359            :out std_logic;
     out360            :out std_logic;
     out361            :out std_logic;
     out362            :out std_logic;
     out363            :out std_logic;
     out364            :out std_logic;
     out365            :out std_logic;
     out366            :out std_logic;
     out367            :out std_logic;
     out368            :out std_logic;
     out369            :out std_logic;
     out370            :out std_logic;
     out371            :out std_logic;
     out372            :out std_logic;
     out373            :out std_logic;
     out374            :out std_logic;
     out375            :out std_logic;
     out376            :out std_logic;
     out377            :out std_logic;
     out378            :out std_logic;
     out379            :out std_logic;
     out380            :out std_logic;
     out381            :out std_logic;
     out382            :out std_logic;
     out383            :out std_logic;
     out384            :out std_logic;
     out385            :out std_logic;
     out386            :out std_logic;
     out387            :out std_logic;
     out388            :out std_logic;
     out389            :out std_logic;
     out390            :out std_logic;
     out391            :out std_logic;
     out392            :out std_logic;
     out393            :out std_logic;
     out394            :out std_logic;
     out395            :out std_logic;
     out396            :out std_logic;
     out397            :out std_logic;
     out398            :out std_logic;
     out399            :out std_logic;
     out400            :out std_logic;
     out401            :out std_logic;
     out402            :out std_logic;
     out403            :out std_logic;
     out404            :out std_logic;
     out405            :out std_logic;
     out406            :out std_logic;
     out407            :out std_logic;
     out408            :out std_logic;
     out409            :out std_logic;
     out410            :out std_logic;
     out411            :out std_logic;
     out412            :out std_logic;
     out413            :out std_logic;
     out414            :out std_logic;
     out415            :out std_logic;
     out416            :out std_logic;
     out417            :out std_logic;
     out418            :out std_logic;
     out419            :out std_logic;
     out420            :out std_logic;
     out421            :out std_logic;
     out422            :out std_logic;
     out423            :out std_logic;
     out424            :out std_logic;
     out425            :out std_logic;
     out426            :out std_logic;
     out427            :out std_logic;
     out428            :out std_logic;
     out429            :out std_logic;
     out430            :out std_logic;
     out431            :out std_logic;
     out432            :out std_logic;
     out433            :out std_logic;
     out434            :out std_logic;
     out435            :out std_logic;
     out436            :out std_logic;
     out437            :out std_logic;
     out438            :out std_logic;
     out439            :out std_logic;
     out440            :out std_logic;
     out441            :out std_logic;
     out442            :out std_logic;
     out443            :out std_logic;
     out444            :out std_logic;
     out445            :out std_logic;
     out446            :out std_logic;
     out447            :out std_logic;
     out448            :out std_logic;
     out449            :out std_logic;
     out450            :out std_logic;
     out451            :out std_logic;
     out452            :out std_logic;
     out453            :out std_logic;
     out454            :out std_logic;
     out455            :out std_logic;
     out456            :out std_logic;
     out457            :out std_logic;
     out458            :out std_logic;
     out459            :out std_logic;
     out460            :out std_logic;
     out461            :out std_logic;
     out462            :out std_logic;
     out463            :out std_logic;
     out464            :out std_logic;
     out465            :out std_logic;
     out466            :out std_logic;
     out467            :out std_logic;
     out468            :out std_logic;
     out469            :out std_logic;
     out470            :out std_logic;
     out471            :out std_logic;
     out472            :out std_logic;
     out473            :out std_logic;
     out474            :out std_logic;
     out475            :out std_logic;
     out476            :out std_logic;
     out477            :out std_logic;
     out478            :out std_logic;
     out479            :out std_logic;
     out480            :out std_logic;
     out481            :out std_logic;
     out482            :out std_logic;
     out483            :out std_logic;
     out484            :out std_logic;
     out485            :out std_logic;
     out486            :out std_logic;
     out487            :out std_logic;
     out488            :out std_logic;
     out489            :out std_logic;
     out490            :out std_logic;
     out491            :out std_logic;
     out492            :out std_logic;
     out493            :out std_logic;
     out494            :out std_logic;
     out495            :out std_logic;
     out496            :out std_logic;
     out497            :out std_logic;
     out498            :out std_logic;
     out499            :out std_logic;
     out500            :out std_logic;
     out501            :out std_logic;
     out502            :out std_logic;
     out503            :out std_logic;
     out504            :out std_logic;
     out505            :out std_logic;
     out506            :out std_logic;
     out507            :out std_logic;
     out508            :out std_logic;
     out509            :out std_logic;
     out510            :out std_logic;
     out511            :out std_logic;
     out512            :out std_logic;
     out513            :out std_logic;
     out514            :out std_logic;
     out515            :out std_logic;
     out516            :out std_logic;
     out517            :out std_logic;
     out518            :out std_logic;
     out519            :out std_logic;
     out520            :out std_logic;
     out521            :out std_logic;
     out522            :out std_logic;
     out523            :out std_logic;
     out524            :out std_logic;
     out525            :out std_logic;
     out526            :out std_logic;
     out527            :out std_logic;
     out528            :out std_logic;
     out529            :out std_logic;
     out530            :out std_logic;
     out531            :out std_logic;
     out532            :out std_logic;
     out533            :out std_logic;
     out534            :out std_logic;
     out535            :out std_logic;
     out536            :out std_logic;
     out537            :out std_logic;
     out538            :out std_logic;
     out539            :out std_logic;
     out540            :out std_logic;
     out541            :out std_logic;
     out542            :out std_logic;
     out543            :out std_logic;
     out544            :out std_logic;
     out545            :out std_logic;
     out546            :out std_logic;
     out547            :out std_logic;
     out548            :out std_logic;
     out549            :out std_logic;
     out550            :out std_logic;
     out551            :out std_logic;
     out552            :out std_logic;
     out553            :out std_logic;
     out554            :out std_logic;
     out555            :out std_logic;
     out556            :out std_logic;
     out557            :out std_logic;
     out558            :out std_logic;
     out559            :out std_logic;
     out560            :out std_logic;
     out561            :out std_logic;
     out562            :out std_logic;
     out563            :out std_logic;
     out564            :out std_logic;
     out565            :out std_logic;
     out566            :out std_logic;
     out567            :out std_logic;
     out568            :out std_logic;
     out569            :out std_logic;
     out570            :out std_logic;
     out571            :out std_logic;
     out572            :out std_logic;
     out573            :out std_logic;
     out574            :out std_logic;
     out575            :out std_logic;
     out576            :out std_logic;
     out577            :out std_logic;
     out578            :out std_logic;
     out579            :out std_logic;
     out580            :out std_logic;
     out581            :out std_logic;
     out582            :out std_logic;
     out583            :out std_logic;
     out584            :out std_logic;
     out585            :out std_logic;
     out586            :out std_logic;
     out587            :out std_logic;
     out588            :out std_logic;
     out589            :out std_logic;
     out590            :out std_logic;
     out591            :out std_logic;
     out592            :out std_logic;
     out593            :out std_logic;
     out594            :out std_logic;
     out595            :out std_logic;
     out596            :out std_logic;
     out597            :out std_logic;
     out598            :out std_logic;
     out599            :out std_logic;
     out600            :out std_logic;
     out601            :out std_logic;
     out602            :out std_logic;
     out603            :out std_logic;
     out604            :out std_logic;
     out605            :out std_logic;
     out606            :out std_logic;
     out607            :out std_logic;
     out608            :out std_logic;
     out609            :out std_logic;
     out610            :out std_logic;
     out611            :out std_logic;
     out612            :out std_logic;
     out613            :out std_logic;
     out614            :out std_logic;
     out615            :out std_logic;
     out616            :out std_logic;
     out617            :out std_logic;
     out618            :out std_logic;
     out619            :out std_logic;
     out620            :out std_logic;
     out621            :out std_logic;
     out622            :out std_logic;
     out623            :out std_logic;
     out624            :out std_logic;
     out625            :out std_logic;
     out626            :out std_logic;
     out627            :out std_logic;
     out628            :out std_logic;
     out629            :out std_logic;
     out630            :out std_logic;
     out631            :out std_logic;
     out632            :out std_logic;
     out633            :out std_logic;
     out634            :out std_logic;
     out635            :out std_logic;
     out636            :out std_logic;
     out637            :out std_logic;
     out638            :out std_logic;
     out639            :out std_logic;
     out640            :out std_logic;
     out641            :out std_logic;
     out642            :out std_logic;
     out643            :out std_logic;
     out644            :out std_logic;
     out645            :out std_logic;
     out646            :out std_logic;
     out647            :out std_logic;
     out648            :out std_logic;
     out649            :out std_logic;
     out650            :out std_logic;
     out651            :out std_logic;
     out652            :out std_logic;
     out653            :out std_logic;
     out654            :out std_logic;
     out655            :out std_logic;
     out656            :out std_logic;
     out657            :out std_logic;
     out658            :out std_logic;
     out659            :out std_logic;
     out660            :out std_logic;
     out661            :out std_logic;
     out662            :out std_logic;
     out663            :out std_logic;
     out664            :out std_logic;
     out665            :out std_logic;
     out666            :out std_logic;
     out667            :out std_logic;
     out668            :out std_logic;
     out669            :out std_logic;
     out670            :out std_logic;
     out671            :out std_logic;
     out672            :out std_logic;
     out673            :out std_logic;
     out674            :out std_logic;
     out675            :out std_logic;
     out676            :out std_logic;
     out677            :out std_logic;
     out678            :out std_logic;
     out679            :out std_logic;
     out680            :out std_logic;
     out681            :out std_logic;
     out682            :out std_logic;
     out683            :out std_logic;
     out684            :out std_logic;
     out685            :out std_logic;
     out686            :out std_logic;
     out687            :out std_logic;
     out688            :out std_logic;
     out689            :out std_logic;
     out690            :out std_logic;
     out691            :out std_logic;
     out692            :out std_logic;
     out693            :out std_logic;
     out694            :out std_logic;
     out695            :out std_logic;
     out696            :out std_logic;
     out697            :out std_logic;
     out698            :out std_logic;
     out699            :out std_logic;
     out700            :out std_logic;
     out701            :out std_logic;
     out702            :out std_logic;
     out703            :out std_logic;
     out704            :out std_logic;
     out705            :out std_logic;
     out706            :out std_logic;
     out707            :out std_logic;
     out708            :out std_logic;
     out709            :out std_logic;
     out710            :out std_logic;
     out711            :out std_logic;
     out712            :out std_logic;
     out713            :out std_logic;
     out714            :out std_logic;
     out715            :out std_logic;
     out716            :out std_logic;
     out717            :out std_logic;
     out718            :out std_logic;
     out719            :out std_logic;
     out720            :out std_logic;
     out721            :out std_logic;
     out722            :out std_logic;
     out723            :out std_logic;
     out724            :out std_logic;
     out725            :out std_logic;
     out726            :out std_logic;
     out727            :out std_logic;
     out728            :out std_logic;
     out729            :out std_logic;
     out730            :out std_logic;
     out731            :out std_logic;
     out732            :out std_logic;
     out733            :out std_logic;
     out734            :out std_logic;
     out735            :out std_logic;
     out736            :out std_logic;
     out737            :out std_logic;
     out738            :out std_logic;
     out739            :out std_logic;
     out740            :out std_logic;
     out741            :out std_logic;
     out742            :out std_logic;
     out743            :out std_logic;
     out744            :out std_logic;
     out745            :out std_logic;
     out746            :out std_logic;
     out747            :out std_logic;
     out748            :out std_logic;
     out749            :out std_logic;
     out750            :out std_logic;
     out751            :out std_logic;
     out752            :out std_logic;
     out753            :out std_logic;
     out754            :out std_logic;
     out755            :out std_logic;
     out756            :out std_logic;
     out757            :out std_logic;
     out758            :out std_logic;
     out759            :out std_logic;
     out760            :out std_logic;
     out761            :out std_logic;
     out762            :out std_logic;
     out763            :out std_logic;
     out764            :out std_logic;
     out765            :out std_logic;
     out766            :out std_logic;
     out767            :out std_logic;
     out768            :out std_logic;
     out769            :out std_logic;
     out770            :out std_logic;
     out771            :out std_logic;
     out772            :out std_logic;
     out773            :out std_logic;
     out774            :out std_logic;
     out775            :out std_logic;
     out776            :out std_logic;
     out777            :out std_logic;
     out778            :out std_logic;
     out779            :out std_logic;
     out780            :out std_logic;
     out781            :out std_logic;
     out782            :out std_logic;
     out783            :out std_logic;
     out784            :out std_logic;
     out785            :out std_logic;
     out786            :out std_logic;
     out787            :out std_logic;
     out788            :out std_logic;
     out789            :out std_logic;
     out790            :out std_logic;
     out791            :out std_logic;
     out792            :out std_logic;
     out793            :out std_logic;
     out794            :out std_logic;
     out795            :out std_logic;
     out796            :out std_logic;
     out797            :out std_logic;
     out798            :out std_logic;
     out799            :out std_logic;
     out800            :out std_logic;
     out801            :out std_logic;
     out802            :out std_logic;
     out803            :out std_logic;
     out804            :out std_logic;
     out805            :out std_logic;
     out806            :out std_logic;
     out807            :out std_logic;
     out808            :out std_logic;
     out809            :out std_logic;
     out810            :out std_logic;
     out811            :out std_logic;
     out812            :out std_logic;
     out813            :out std_logic;
     out814            :out std_logic;
     out815            :out std_logic;
     out816            :out std_logic;
     out817            :out std_logic;
     out818            :out std_logic;
     out819            :out std_logic;
     out820            :out std_logic;
     out821            :out std_logic;
     out822            :out std_logic;
     out823            :out std_logic;
     out824            :out std_logic;
     out825            :out std_logic;
     out826            :out std_logic;
     out827            :out std_logic;
     out828            :out std_logic;
     out829            :out std_logic;
     out830            :out std_logic;
     out831            :out std_logic;
     out832            :out std_logic;
     out833            :out std_logic;
     out834            :out std_logic;
     out835            :out std_logic;
     out836            :out std_logic;
     out837            :out std_logic;
     out838            :out std_logic;
     out839            :out std_logic;
     out840            :out std_logic;
     out841            :out std_logic;
     out842            :out std_logic;
     out843            :out std_logic;
     out844            :out std_logic;
     out845            :out std_logic;
     out846            :out std_logic;
     out847            :out std_logic;
     out848            :out std_logic;
     out849            :out std_logic;
     out850            :out std_logic;
     out851            :out std_logic;
     out852            :out std_logic;
     out853            :out std_logic;
     out854            :out std_logic;
     out855            :out std_logic;
     out856            :out std_logic;
     out857            :out std_logic;
     out858            :out std_logic;
     out859            :out std_logic;
     out860            :out std_logic;
     out861            :out std_logic;
     out862            :out std_logic;
     out863            :out std_logic;
     out864            :out std_logic;
     out865            :out std_logic;
     out866            :out std_logic;
     out867            :out std_logic;
     out868            :out std_logic;
     out869            :out std_logic;
     out870            :out std_logic;
     out871            :out std_logic;
     out872            :out std_logic;
     out873            :out std_logic;
     out874            :out std_logic;
     out875            :out std_logic;
     out876            :out std_logic;
     out877            :out std_logic;
     out878            :out std_logic;
     out879            :out std_logic;
     out880            :out std_logic;
     out881            :out std_logic;
     out882            :out std_logic;
     out883            :out std_logic;
     out884            :out std_logic;
     out885            :out std_logic;
     out886            :out std_logic;
     out887            :out std_logic;
     out888            :out std_logic;
     out889            :out std_logic;
     out890            :out std_logic;
     out891            :out std_logic;
     out892            :out std_logic;
     out893            :out std_logic;
     out894            :out std_logic;
     out895            :out std_logic;
     out896            :out std_logic;
     out897            :out std_logic;
     out898            :out std_logic;
     out899            :out std_logic;
     out900            :out std_logic;
     out901            :out std_logic;
     out902            :out std_logic;
     out903            :out std_logic;
     out904            :out std_logic;
     out905            :out std_logic;
     out906            :out std_logic;
     out907            :out std_logic;
     out908            :out std_logic;
     out909            :out std_logic;
     out910            :out std_logic;
     out911            :out std_logic;
     out912            :out std_logic;
     out913            :out std_logic;
     out914            :out std_logic;
     out915            :out std_logic;
     out916            :out std_logic;
     out917            :out std_logic;
     out918            :out std_logic;
     out919            :out std_logic;
     out920            :out std_logic;
     out921            :out std_logic;
     out922            :out std_logic;
     out923            :out std_logic;
     out924            :out std_logic;
     out925            :out std_logic;
     out926            :out std_logic;
     out927            :out std_logic;
     out928            :out std_logic;
     out929            :out std_logic;
     out930            :out std_logic;
     out931            :out std_logic;
     out932            :out std_logic;
     out933            :out std_logic;
     out934            :out std_logic;
     out935            :out std_logic;
     out936            :out std_logic;
     out937            :out std_logic;
     out938            :out std_logic;
     out939            :out std_logic;
     out940            :out std_logic;
     out941            :out std_logic;
     out942            :out std_logic;
     out943            :out std_logic;
     out944            :out std_logic;
     out945            :out std_logic;
     out946            :out std_logic;
     out947            :out std_logic;
     out948            :out std_logic;
     out949            :out std_logic;
     out950            :out std_logic;
     out951            :out std_logic;
     out952            :out std_logic;
     out953            :out std_logic;
     out954            :out std_logic;
     out955            :out std_logic;
     out956            :out std_logic;
     out957            :out std_logic;
     out958            :out std_logic;
     out959            :out std_logic;
     out960            :out std_logic;
     out961            :out std_logic;
     out962            :out std_logic;
     out963            :out std_logic;
     out964            :out std_logic;
     out965            :out std_logic;
     out966            :out std_logic;
     out967            :out std_logic;
     out968            :out std_logic;
     out969            :out std_logic;
     out970            :out std_logic;
     out971            :out std_logic;
     out972            :out std_logic;
     out973            :out std_logic;
     out974            :out std_logic;
     out975            :out std_logic;
     out976            :out std_logic;
     out977            :out std_logic;
     out978            :out std_logic;
     out979            :out std_logic;
     out980            :out std_logic;
     out981            :out std_logic;
     out982            :out std_logic;
     out983            :out std_logic;
     out984            :out std_logic;
     out985            :out std_logic;
     out986            :out std_logic;
     out987            :out std_logic;
     out988            :out std_logic;
     out989            :out std_logic;
     out990            :out std_logic;
     out991            :out std_logic;
     out992            :out std_logic;
     out993            :out std_logic;
     out994            :out std_logic;
     out995            :out std_logic;
     out996            :out std_logic;
     out997            :out std_logic;
     out998            :out std_logic;
     out999            :out std_logic;
     out1000            :out std_logic;
     out1001            :out std_logic;
     out1002            :out std_logic;
     out1003            :out std_logic;
     out1004            :out std_logic;
     out1005            :out std_logic;
     out1006            :out std_logic;
     out1007            :out std_logic;
     out1008            :out std_logic;
     out1009            :out std_logic;
     out1010            :out std_logic;
     out1011            :out std_logic;
     out1012            :out std_logic;
     out1013            :out std_logic;
     out1014            :out std_logic;
     out1015            :out std_logic;
     out1016            :out std_logic;
     out1017            :out std_logic;
     out1018            :out std_logic;
     out1019            :out std_logic;
     out1020            :out std_logic;
     out1021            :out std_logic;
     out1022            :out std_logic;
     out1023            :out std_logic;
     out1024            :out std_logic;
     out1025            :out std_logic;
     out1026            :out std_logic;
     out1027            :out std_logic;
     out1028            :out std_logic;
     out1029            :out std_logic;
     out1030            :out std_logic;
     out1031            :out std_logic;
     out1032            :out std_logic;
     out1033            :out std_logic;
     out1034            :out std_logic;
     out1035            :out std_logic;
     out1036            :out std_logic;
     out1037            :out std_logic;
     out1038            :out std_logic;
     out1039            :out std_logic;
     out1040            :out std_logic;
     out1041            :out std_logic;
     out1042            :out std_logic;
     out1043            :out std_logic;
     out1044            :out std_logic;
     out1045            :out std_logic;
     out1046            :out std_logic;
     out1047            :out std_logic;
     out1048            :out std_logic;
     out1049            :out std_logic;
     out1050            :out std_logic;
     out1051            :out std_logic;
     out1052            :out std_logic;
     out1053            :out std_logic;
     out1054            :out std_logic;
     out1055            :out std_logic;
     out1056            :out std_logic;
     out1057            :out std_logic;
     out1058            :out std_logic;
     out1059            :out std_logic;
     out1060            :out std_logic;
     out1061            :out std_logic;
     out1062            :out std_logic;
     out1063            :out std_logic;
     out1064            :out std_logic;
     out1065            :out std_logic;
     out1066            :out std_logic;
     out1067            :out std_logic;
     out1068            :out std_logic;
     out1069            :out std_logic;
     out1070            :out std_logic;
     out1071            :out std_logic;
     out1072            :out std_logic;
     out1073            :out std_logic;
     out1074            :out std_logic;
     out1075            :out std_logic;
     out1076            :out std_logic;
     out1077            :out std_logic;
     out1078            :out std_logic;
     out1079            :out std_logic;
     out1080            :out std_logic;
     out1081            :out std_logic;
     out1082            :out std_logic;
     out1083            :out std_logic;
     out1084            :out std_logic;
     out1085            :out std_logic;
     out1086            :out std_logic;
     out1087            :out std_logic;
     out1088            :out std_logic;
     out1089            :out std_logic;
     out1090            :out std_logic;
     out1091            :out std_logic;
     out1092            :out std_logic;
     out1093            :out std_logic;
     out1094            :out std_logic;
     out1095            :out std_logic;
     out1096            :out std_logic;
     out1097            :out std_logic;
     out1098            :out std_logic;
     out1099            :out std_logic;
     out1100            :out std_logic;
     out1101            :out std_logic;
     out1102            :out std_logic;
     out1103            :out std_logic;
     out1104            :out std_logic;
     out1105            :out std_logic;
     out1106            :out std_logic;
     out1107            :out std_logic;
     out1108            :out std_logic;
     out1109            :out std_logic;
     out1110            :out std_logic;
     out1111            :out std_logic;
     out1112            :out std_logic;
     out1113            :out std_logic;
     out1114            :out std_logic;
     out1115            :out std_logic;
     out1116            :out std_logic;
     out1117            :out std_logic;
     out1118            :out std_logic;
     out1119            :out std_logic;
     out1120            :out std_logic;
     out1121            :out std_logic;
     out1122            :out std_logic;
     out1123            :out std_logic;
     out1124            :out std_logic;
     out1125            :out std_logic;
     out1126            :out std_logic;
     out1127            :out std_logic;
     out1128            :out std_logic;
     out1129            :out std_logic;
     out1130            :out std_logic;
     out1131            :out std_logic;
     out1132            :out std_logic;
     out1133            :out std_logic;
     out1134            :out std_logic;
     out1135            :out std_logic;
     out1136            :out std_logic;
     out1137            :out std_logic;
     out1138            :out std_logic;
     out1139            :out std_logic;
     out1140            :out std_logic;
     out1141            :out std_logic;
     out1142            :out std_logic;
     out1143            :out std_logic;
     out1144            :out std_logic;
     out1145            :out std_logic;
     out1146            :out std_logic;
     out1147            :out std_logic;
     out1148            :out std_logic;
     out1149            :out std_logic;
     out1150            :out std_logic;
     out1151            :out std_logic;
     out1152            :out std_logic;
     out1153            :out std_logic;
     out1154            :out std_logic;
     out1155            :out std_logic;
     out1156            :out std_logic;
     out1157            :out std_logic;
     out1158            :out std_logic;
     out1159            :out std_logic;
     out1160            :out std_logic;
     out1161            :out std_logic;
     out1162            :out std_logic;
     out1163            :out std_logic;
     out1164            :out std_logic;
     out1165            :out std_logic;
     out1166            :out std_logic;
     out1167            :out std_logic;
     out1168            :out std_logic;
     out1169            :out std_logic;
     out1170            :out std_logic;
     out1171            :out std_logic;
     out1172            :out std_logic;
     out1173            :out std_logic;
     out1174            :out std_logic;
     out1175            :out std_logic;
     out1176            :out std_logic;
     out1177            :out std_logic;
     out1178            :out std_logic;
     out1179            :out std_logic;
     out1180            :out std_logic;
     out1181            :out std_logic;
     out1182            :out std_logic;
     out1183            :out std_logic;
     out1184            :out std_logic;
     out1185            :out std_logic;
     out1186            :out std_logic;
     out1187            :out std_logic;
     out1188            :out std_logic;
     out1189            :out std_logic;
     out1190            :out std_logic;
     out1191            :out std_logic;
     out1192            :out std_logic;
     out1193            :out std_logic;
     out1194            :out std_logic;
     out1195            :out std_logic;
     out1196            :out std_logic;
     out1197            :out std_logic;
     out1198            :out std_logic;
     out1199            :out std_logic;
     out1200            :out std_logic;
     out1201            :out std_logic;
     out1202            :out std_logic;
     out1203            :out std_logic;
     out1204            :out std_logic;
     out1205            :out std_logic;
     out1206            :out std_logic;
     out1207            :out std_logic;
     out1208            :out std_logic;
     out1209            :out std_logic;
     out1210            :out std_logic;
     out1211            :out std_logic;
     out1212            :out std_logic;
     out1213            :out std_logic;
     out1214            :out std_logic;
     out1215            :out std_logic;
     out1216            :out std_logic;
     out1217            :out std_logic;
     out1218            :out std_logic;
     out1219            :out std_logic;
     out1220            :out std_logic;
     out1221            :out std_logic;
     out1222            :out std_logic;
     out1223            :out std_logic;
     out1224            :out std_logic;
     out1225            :out std_logic;
     out1226            :out std_logic;
     out1227            :out std_logic;
     out1228            :out std_logic;
     out1229            :out std_logic;
     out1230            :out std_logic;
     out1231            :out std_logic;
     out1232            :out std_logic;
     out1233            :out std_logic;
     out1234            :out std_logic;
     out1235            :out std_logic;
     out1236            :out std_logic;
     out1237            :out std_logic;
     out1238            :out std_logic;
     out1239            :out std_logic;
     out1240            :out std_logic;
     out1241            :out std_logic;
     out1242            :out std_logic;
     out1243            :out std_logic;
     out1244            :out std_logic;
     out1245            :out std_logic;
     out1246            :out std_logic;
     out1247            :out std_logic;
     out1248            :out std_logic;
     out1249            :out std_logic;
     out1250            :out std_logic;
     out1251            :out std_logic;
     out1252            :out std_logic;
     out1253            :out std_logic;
     out1254            :out std_logic;
     out1255            :out std_logic;
     out1256            :out std_logic;
     out1257            :out std_logic;
     out1258            :out std_logic;
     out1259            :out std_logic;
     out1260            :out std_logic;
     out1261            :out std_logic;
     out1262            :out std_logic;
     out1263            :out std_logic;
     out1264            :out std_logic;
     out1265            :out std_logic;
     out1266            :out std_logic;
     out1267            :out std_logic;
     out1268            :out std_logic;
     out1269            :out std_logic;
     out1270            :out std_logic;
     out1271            :out std_logic;
     out1272            :out std_logic;
     out1273            :out std_logic;
     out1274            :out std_logic;
     out1275            :out std_logic;
     out1276            :out std_logic;
     out1277            :out std_logic;
     out1278            :out std_logic;
     out1279            :out std_logic;
     out1280            :out std_logic;
     out1281            :out std_logic;
     out1282            :out std_logic;
     out1283            :out std_logic;
     out1284            :out std_logic;
     out1285            :out std_logic;
     out1286            :out std_logic;
     out1287            :out std_logic;
     out1288            :out std_logic;
     out1289            :out std_logic;
     out1290            :out std_logic;
     out1291            :out std_logic;
     out1292            :out std_logic;
     out1293            :out std_logic;
     out1294            :out std_logic;
     out1295            :out std_logic;
     out1296            :out std_logic;
     out1297            :out std_logic;
     out1298            :out std_logic;
     out1299            :out std_logic;
     out1300            :out std_logic;
     out1301            :out std_logic;
     out1302            :out std_logic;
     out1303            :out std_logic;
     out1304            :out std_logic;
     out1305            :out std_logic;
     out1306            :out std_logic;
     out1307            :out std_logic;
     out1308            :out std_logic;
     out1309            :out std_logic;
     out1310            :out std_logic;
     out1311            :out std_logic;
     out1312            :out std_logic;
     out1313            :out std_logic;
     out1314            :out std_logic;
     out1315            :out std_logic;
     out1316            :out std_logic;
     out1317            :out std_logic;
     out1318            :out std_logic;
     out1319            :out std_logic;
     out1320            :out std_logic;
     out1321            :out std_logic;
     out1322            :out std_logic;
     out1323            :out std_logic;
     out1324            :out std_logic;
     out1325            :out std_logic;
     out1326            :out std_logic;
     out1327            :out std_logic;
     out1328            :out std_logic;
     out1329            :out std_logic;
     out1330            :out std_logic;
     out1331            :out std_logic;
     out1332            :out std_logic;
     out1333            :out std_logic;
     out1334            :out std_logic;
     out1335            :out std_logic;
     out1336            :out std_logic;
     out1337            :out std_logic;
     out1338            :out std_logic;
     out1339            :out std_logic;
     out1340            :out std_logic;
     out1341            :out std_logic;
     out1342            :out std_logic;
     out1343            :out std_logic;
     out1344            :out std_logic;
     out1345            :out std_logic;
     out1346            :out std_logic;
     out1347            :out std_logic;
     out1348            :out std_logic;
     out1349            :out std_logic;
     out1350            :out std_logic;
     out1351            :out std_logic;
     out1352            :out std_logic;
     out1353            :out std_logic;
     out1354            :out std_logic;
     out1355            :out std_logic;
     out1356            :out std_logic;
     out1357            :out std_logic;
     out1358            :out std_logic;
     out1359            :out std_logic;
     out1360            :out std_logic;
     out1361            :out std_logic;
     out1362            :out std_logic;
     out1363            :out std_logic;
     out1364            :out std_logic;
     out1365            :out std_logic;
     out1366            :out std_logic;
     out1367            :out std_logic;
     out1368            :out std_logic;
     out1369            :out std_logic;
     out1370            :out std_logic;
     out1371            :out std_logic;
     out1372            :out std_logic;
     out1373            :out std_logic;
     out1374            :out std_logic;
     out1375            :out std_logic;
     out1376            :out std_logic;
     out1377            :out std_logic;
     out1378            :out std_logic;
     out1379            :out std_logic;
     out1380            :out std_logic;
     out1381            :out std_logic;
     out1382            :out std_logic;
     out1383            :out std_logic;
     out1384            :out std_logic;
     out1385            :out std_logic;
     out1386            :out std_logic;
     out1387            :out std_logic;
     out1388            :out std_logic;
     out1389            :out std_logic;
     out1390            :out std_logic;
     out1391            :out std_logic;
     out1392            :out std_logic;
     out1393            :out std_logic;
     out1394            :out std_logic;
     out1395            :out std_logic;
     out1396            :out std_logic;
     out1397            :out std_logic;
     out1398            :out std_logic;
     out1399            :out std_logic;
     out1400            :out std_logic;
     out1401            :out std_logic;
     out1402            :out std_logic;
     out1403            :out std_logic;
     out1404            :out std_logic;
     out1405            :out std_logic;
     out1406            :out std_logic;
     out1407            :out std_logic;
     out1408            :out std_logic;
     out1409            :out std_logic;
     out1410            :out std_logic;
     out1411            :out std_logic;
     out1412            :out std_logic;
     out1413            :out std_logic;
     out1414            :out std_logic;
     out1415            :out std_logic;
     out1416            :out std_logic;
     out1417            :out std_logic;
     out1418            :out std_logic;
     out1419            :out std_logic;
     out1420            :out std_logic;
     out1421            :out std_logic;
     out1422            :out std_logic;
     out1423            :out std_logic;
     out1424            :out std_logic;
     out1425            :out std_logic;
     out1426            :out std_logic;
     out1427            :out std_logic;
     out1428            :out std_logic;
     out1429            :out std_logic;
     out1430            :out std_logic;
     out1431            :out std_logic;
     out1432            :out std_logic;
     out1433            :out std_logic;
     out1434            :out std_logic;
     out1435            :out std_logic;
     out1436            :out std_logic;
     out1437            :out std_logic;
     out1438            :out std_logic;
     out1439            :out std_logic;
     out1440            :out std_logic;
     out1441            :out std_logic;
     out1442            :out std_logic;
     out1443            :out std_logic;
     out1444            :out std_logic;
     out1445            :out std_logic;
     out1446            :out std_logic;
     out1447            :out std_logic;
     out1448            :out std_logic;
     out1449            :out std_logic;
     out1450            :out std_logic;
     out1451            :out std_logic;
     out1452            :out std_logic;
     out1453            :out std_logic;
     out1454            :out std_logic;
     out1455            :out std_logic;
     out1456            :out std_logic;
     out1457            :out std_logic;
     out1458            :out std_logic;
     out1459            :out std_logic;
     out1460            :out std_logic;
     out1461            :out std_logic;
     out1462            :out std_logic;
     out1463            :out std_logic;
     out1464            :out std_logic;
     out1465            :out std_logic;
     out1466            :out std_logic;
     out1467            :out std_logic;
     out1468            :out std_logic;
     out1469            :out std_logic;
     out1470            :out std_logic;
     out1471            :out std_logic;
     out1472            :out std_logic;
     out1473            :out std_logic;
     out1474            :out std_logic;
     out1475            :out std_logic;
     out1476            :out std_logic;
     out1477            :out std_logic;
     out1478            :out std_logic;
     out1479            :out std_logic;
     out1480            :out std_logic;
     out1481            :out std_logic;
     out1482            :out std_logic;
     out1483            :out std_logic;
     out1484            :out std_logic;
     out1485            :out std_logic;
     out1486            :out std_logic;
     out1487            :out std_logic;
     out1488            :out std_logic;
     out1489            :out std_logic;
     out1490            :out std_logic;
     out1491            :out std_logic;
     out1492            :out std_logic;
     out1493            :out std_logic;
     out1494            :out std_logic;
     out1495            :out std_logic;
     out1496            :out std_logic;
     out1497            :out std_logic;
     out1498            :out std_logic;
     out1499            :out std_logic;
     out1500            :out std_logic;
     out1501            :out std_logic;
     out1502            :out std_logic;
     out1503            :out std_logic;
     out1504            :out std_logic;
     out1505            :out std_logic;
     out1506            :out std_logic;
     out1507            :out std_logic;
     out1508            :out std_logic;
     out1509            :out std_logic;
     out1510            :out std_logic;
     out1511            :out std_logic;
     out1512            :out std_logic;
     out1513            :out std_logic;
     out1514            :out std_logic;
     out1515            :out std_logic;
     out1516            :out std_logic;
     out1517            :out std_logic;
     out1518            :out std_logic;
     out1519            :out std_logic;
     out1520            :out std_logic;
     out1521            :out std_logic;
     out1522            :out std_logic;
     out1523            :out std_logic;
     out1524            :out std_logic;
     out1525            :out std_logic;
     out1526            :out std_logic;
     out1527            :out std_logic;
     out1528            :out std_logic;
     out1529            :out std_logic;
     out1530            :out std_logic;
     out1531            :out std_logic;
     out1532            :out std_logic;
     out1533            :out std_logic;
     out1534            :out std_logic;
     out1535            :out std_logic;
     out1536            :out std_logic;
     out1537            :out std_logic;
     out1538            :out std_logic;
     out1539            :out std_logic;
     out1540            :out std_logic;
     out1541            :out std_logic;
     out1542            :out std_logic;
     out1543            :out std_logic;
     out1544            :out std_logic;
     out1545            :out std_logic;
     out1546            :out std_logic;
     out1547            :out std_logic;
     out1548            :out std_logic;
     out1549            :out std_logic;
     out1550            :out std_logic;
     out1551            :out std_logic;
     out1552            :out std_logic;
     out1553            :out std_logic;
     out1554            :out std_logic;
     out1555            :out std_logic;
     out1556            :out std_logic;
     out1557            :out std_logic;
     out1558            :out std_logic;
     out1559            :out std_logic;
     out1560            :out std_logic;
     out1561            :out std_logic;
     out1562            :out std_logic;
     out1563            :out std_logic;
     out1564            :out std_logic;
     out1565            :out std_logic;
     out1566            :out std_logic;
     out1567            :out std_logic;
     out1568            :out std_logic;
     out1569            :out std_logic;
     out1570            :out std_logic;
     out1571            :out std_logic;
     out1572            :out std_logic;
     out1573            :out std_logic;
     out1574            :out std_logic;
     out1575            :out std_logic;
     out1576            :out std_logic;
     out1577            :out std_logic;
     out1578            :out std_logic;
     out1579            :out std_logic;
     out1580            :out std_logic;
     out1581            :out std_logic;
     out1582            :out std_logic;
     out1583            :out std_logic;
     out1584            :out std_logic;
     out1585            :out std_logic;
     out1586            :out std_logic;
     out1587            :out std_logic;
     out1588            :out std_logic;
     out1589            :out std_logic;
     out1590            :out std_logic;
     out1591            :out std_logic;
     out1592            :out std_logic;
     out1593            :out std_logic;
     out1594            :out std_logic;
     out1595            :out std_logic;
     out1596            :out std_logic;
     out1597            :out std_logic;
     out1598            :out std_logic;
     out1599            :out std_logic;
     out1600            :out std_logic;
     out1601            :out std_logic;
     out1602            :out std_logic;
     out1603            :out std_logic;
     out1604            :out std_logic;
     out1605            :out std_logic;
     out1606            :out std_logic;
     out1607            :out std_logic;
     out1608            :out std_logic;
     out1609            :out std_logic;
     out1610            :out std_logic;
     out1611            :out std_logic;
     out1612            :out std_logic;
     out1613            :out std_logic;
     out1614            :out std_logic;
     out1615            :out std_logic;
     out1616            :out std_logic;
     out1617            :out std_logic;
     out1618            :out std_logic;
     out1619            :out std_logic;
     out1620            :out std_logic;
     out1621            :out std_logic;
     out1622            :out std_logic;
     out1623            :out std_logic;
     out1624            :out std_logic;
     out1625            :out std_logic;
     out1626            :out std_logic;
     out1627            :out std_logic;
     out1628            :out std_logic;
     out1629            :out std_logic;
     out1630            :out std_logic;
     out1631            :out std_logic;
     out1632            :out std_logic;
     out1633            :out std_logic;
     out1634            :out std_logic;
     out1635            :out std_logic;
     out1636            :out std_logic;
     out1637            :out std_logic;
     out1638            :out std_logic;
     out1639            :out std_logic;
     out1640            :out std_logic;
     out1641            :out std_logic;
     out1642            :out std_logic;
     out1643            :out std_logic;
     out1644            :out std_logic;
     out1645            :out std_logic;
     out1646            :out std_logic;
     out1647            :out std_logic;
     out1648            :out std_logic;
     out1649            :out std_logic;
     out1650            :out std_logic;
     out1651            :out std_logic;
     out1652            :out std_logic;
     out1653            :out std_logic;
     out1654            :out std_logic;
     out1655            :out std_logic;
     out1656            :out std_logic;
     out1657            :out std_logic;
     out1658            :out std_logic;
     out1659            :out std_logic;
     out1660            :out std_logic;
     out1661            :out std_logic;
     out1662            :out std_logic;
     out1663            :out std_logic;
     out1664            :out std_logic;
     out1665            :out std_logic;
     out1666            :out std_logic;
     out1667            :out std_logic;
     out1668            :out std_logic;
     out1669            :out std_logic;
     out1670            :out std_logic;
     out1671            :out std_logic;
     out1672            :out std_logic;
     out1673            :out std_logic;
     out1674            :out std_logic;
     out1675            :out std_logic;
     out1676            :out std_logic;
     out1677            :out std_logic;
     out1678            :out std_logic;
     out1679            :out std_logic;
     out1680            :out std_logic;
     out1681            :out std_logic;
     out1682            :out std_logic;
     out1683            :out std_logic;
     out1684            :out std_logic;
     out1685            :out std_logic;
     out1686            :out std_logic;
     out1687            :out std_logic;
     out1688            :out std_logic;
     out1689            :out std_logic;
     out1690            :out std_logic;
     out1691            :out std_logic;
     out1692            :out std_logic;
     out1693            :out std_logic;
     out1694            :out std_logic;
     out1695            :out std_logic;
     out1696            :out std_logic;
     out1697            :out std_logic;
     out1698            :out std_logic;
     out1699            :out std_logic;
     out1700            :out std_logic;
     out1701            :out std_logic;
     out1702            :out std_logic;
     out1703            :out std_logic;
     out1704            :out std_logic;
     out1705            :out std_logic;
     out1706            :out std_logic;
     out1707            :out std_logic;
     out1708            :out std_logic;
     out1709            :out std_logic;
     out1710            :out std_logic;
     out1711            :out std_logic;
     out1712            :out std_logic;
     out1713            :out std_logic;
     out1714            :out std_logic;
     out1715            :out std_logic;
     out1716            :out std_logic;
     out1717            :out std_logic;
     out1718            :out std_logic;
     out1719            :out std_logic;
     out1720            :out std_logic;
     out1721            :out std_logic;
     out1722            :out std_logic;
     out1723            :out std_logic;
     out1724            :out std_logic;
     out1725            :out std_logic;
     out1726            :out std_logic;
     out1727            :out std_logic;
     out1728            :out std_logic;
     out1729            :out std_logic;
     out1730            :out std_logic;
     out1731            :out std_logic;
     out1732            :out std_logic;
     out1733            :out std_logic;
     out1734            :out std_logic;
     out1735            :out std_logic;
     out1736            :out std_logic;
     out1737            :out std_logic;
     out1738            :out std_logic;
     out1739            :out std_logic;
     out1740            :out std_logic;
     out1741            :out std_logic;
     out1742            :out std_logic;
     out1743            :out std_logic;
     out1744            :out std_logic;
     out1745            :out std_logic;
     out1746            :out std_logic;
     out1747            :out std_logic;
     out1748            :out std_logic;
     out1749            :out std_logic;
     out1750            :out std_logic;
     out1751            :out std_logic;
     out1752            :out std_logic;
     out1753            :out std_logic;
     out1754            :out std_logic;
     out1755            :out std_logic;
     out1756            :out std_logic;
     out1757            :out std_logic;
     out1758            :out std_logic;
     out1759            :out std_logic;
     out1760            :out std_logic;
     out1761            :out std_logic;
     out1762            :out std_logic;
     out1763            :out std_logic;
     out1764            :out std_logic;
     out1765            :out std_logic;
     out1766            :out std_logic;
     out1767            :out std_logic;
     out1768            :out std_logic;
     out1769            :out std_logic;
     out1770            :out std_logic;
     out1771            :out std_logic;
     out1772            :out std_logic;
     out1773            :out std_logic;
     out1774            :out std_logic;
     out1775            :out std_logic;
     out1776            :out std_logic;
     out1777            :out std_logic;
     out1778            :out std_logic;
     out1779            :out std_logic;
     out1780            :out std_logic;
     out1781            :out std_logic;
     out1782            :out std_logic;
     out1783            :out std_logic;
     out1784            :out std_logic;
     out1785            :out std_logic;
     out1786            :out std_logic;
     out1787            :out std_logic;
     out1788            :out std_logic;
     out1789            :out std_logic;
     out1790            :out std_logic;
     out1791            :out std_logic;
     out1792            :out std_logic;
     out1793            :out std_logic;
     out1794            :out std_logic;
     out1795            :out std_logic;
     out1796            :out std_logic;
     out1797            :out std_logic;
     out1798            :out std_logic;
     out1799            :out std_logic;
     out1800            :out std_logic;
     out1801            :out std_logic;
     out1802            :out std_logic;
     out1803            :out std_logic;
     out1804            :out std_logic;
     out1805            :out std_logic;
     out1806            :out std_logic;
     out1807            :out std_logic;
     out1808            :out std_logic;
     out1809            :out std_logic;
     out1810            :out std_logic;
     out1811            :out std_logic;
     out1812            :out std_logic;
     out1813            :out std_logic;
     out1814            :out std_logic;
     out1815            :out std_logic;
     out1816            :out std_logic;
     out1817            :out std_logic;
     out1818            :out std_logic;
     out1819            :out std_logic;
     out1820            :out std_logic;
     out1821            :out std_logic;
     out1822            :out std_logic;
     out1823            :out std_logic;
     out1824            :out std_logic;
     out1825            :out std_logic;
     out1826            :out std_logic;
     out1827            :out std_logic;
     out1828            :out std_logic;
     out1829            :out std_logic;
     out1830            :out std_logic;
     out1831            :out std_logic;
     out1832            :out std_logic;
     out1833            :out std_logic;
     out1834            :out std_logic;
     out1835            :out std_logic;
     out1836            :out std_logic;
     out1837            :out std_logic;
     out1838            :out std_logic;
     out1839            :out std_logic;
     out1840            :out std_logic;
     out1841            :out std_logic;
     out1842            :out std_logic;
     out1843            :out std_logic;
     out1844            :out std_logic;
     out1845            :out std_logic;
     out1846            :out std_logic;
     out1847            :out std_logic;
     out1848            :out std_logic;
     out1849            :out std_logic;
     out1850            :out std_logic;
     out1851            :out std_logic;
     out1852            :out std_logic;
     out1853            :out std_logic;
     out1854            :out std_logic;
     out1855            :out std_logic;
     out1856            :out std_logic;
     out1857            :out std_logic;
     out1858            :out std_logic;
     out1859            :out std_logic;
     out1860            :out std_logic;
     out1861            :out std_logic;
     out1862            :out std_logic;
     out1863            :out std_logic;
     out1864            :out std_logic;
     out1865            :out std_logic;
     out1866            :out std_logic;
     out1867            :out std_logic;
     out1868            :out std_logic;
     out1869            :out std_logic;
     out1870            :out std_logic;
     out1871            :out std_logic;
     out1872            :out std_logic;
     out1873            :out std_logic;
     out1874            :out std_logic;
     out1875            :out std_logic;
     out1876            :out std_logic;
     out1877            :out std_logic;
     out1878            :out std_logic;
     out1879            :out std_logic;
     out1880            :out std_logic;
     out1881            :out std_logic;
     out1882            :out std_logic;
     out1883            :out std_logic;
     out1884            :out std_logic;
     out1885            :out std_logic;
     out1886            :out std_logic;
     out1887            :out std_logic;
     out1888            :out std_logic;
     out1889            :out std_logic;
     out1890            :out std_logic;
     out1891            :out std_logic;
     out1892            :out std_logic;
     out1893            :out std_logic;
     out1894            :out std_logic;
     out1895            :out std_logic;
     out1896            :out std_logic;
     out1897            :out std_logic;
     out1898            :out std_logic;
     out1899            :out std_logic;
     out1900            :out std_logic;
     out1901            :out std_logic;
     out1902            :out std_logic;
     out1903            :out std_logic;
     out1904            :out std_logic;
     out1905            :out std_logic;
     out1906            :out std_logic;
     out1907            :out std_logic;
     out1908            :out std_logic;
     out1909            :out std_logic;
     out1910            :out std_logic;
     out1911            :out std_logic;
     out1912            :out std_logic;
     out1913            :out std_logic;
     out1914            :out std_logic;
     out1915            :out std_logic;
     out1916            :out std_logic;
     out1917            :out std_logic;
     out1918            :out std_logic;
     out1919            :out std_logic;
     out1920            :out std_logic;
     out1921            :out std_logic;
     out1922            :out std_logic;
     out1923            :out std_logic;
     out1924            :out std_logic;
     out1925            :out std_logic;
     out1926            :out std_logic;
     out1927            :out std_logic;
     out1928            :out std_logic;
     out1929            :out std_logic;
     out1930            :out std_logic;
     out1931            :out std_logic;
     out1932            :out std_logic;
     out1933            :out std_logic;
     out1934            :out std_logic;
     out1935            :out std_logic;
     out1936            :out std_logic;
     out1937            :out std_logic;
     out1938            :out std_logic;
     out1939            :out std_logic;
     out1940            :out std_logic;
     out1941            :out std_logic;
     out1942            :out std_logic;
     out1943            :out std_logic;
     out1944            :out std_logic;
     out1945            :out std_logic;
     out1946            :out std_logic;
     out1947            :out std_logic;
     out1948            :out std_logic;
     out1949            :out std_logic;
     out1950            :out std_logic;
     out1951            :out std_logic;
     out1952            :out std_logic;
     out1953            :out std_logic;
     out1954            :out std_logic;
     out1955            :out std_logic;
     out1956            :out std_logic;
     out1957            :out std_logic;
     out1958            :out std_logic;
     out1959            :out std_logic;
     out1960            :out std_logic;
     out1961            :out std_logic;
     out1962            :out std_logic;
     out1963            :out std_logic;
     out1964            :out std_logic;
     out1965            :out std_logic;
     out1966            :out std_logic;
     out1967            :out std_logic;
     out1968            :out std_logic;
     out1969            :out std_logic;
     out1970            :out std_logic;
     out1971            :out std_logic;
     out1972            :out std_logic;
     out1973            :out std_logic;
     out1974            :out std_logic;
     out1975            :out std_logic;
     out1976            :out std_logic;
     out1977            :out std_logic;
     out1978            :out std_logic;
     out1979            :out std_logic;
     out1980            :out std_logic;
     out1981            :out std_logic;
     out1982            :out std_logic;
     out1983            :out std_logic;
     out1984            :out std_logic;
     out1985            :out std_logic;
     out1986            :out std_logic;
     out1987            :out std_logic;
     out1988            :out std_logic;
     out1989            :out std_logic;
     out1990            :out std_logic;
     out1991            :out std_logic;
     out1992            :out std_logic;
     out1993            :out std_logic;
     out1994            :out std_logic;
     out1995            :out std_logic;
     out1996            :out std_logic;
     out1997            :out std_logic;
     out1998            :out std_logic;
     out1999            :out std_logic;
     out2000            :out std_logic;
     out2001            :out std_logic;
     out2002            :out std_logic;
     out2003            :out std_logic;
     out2004            :out std_logic;
     out2005            :out std_logic;
     out2006            :out std_logic;
     out2007            :out std_logic;
     out2008            :out std_logic;
     out2009            :out std_logic;
     out2010            :out std_logic;
     out2011            :out std_logic;
     out2012            :out std_logic;
     out2013            :out std_logic;
     out2014            :out std_logic;
     out2015            :out std_logic;
     out2016            :out std_logic;
     out2017            :out std_logic;
     out2018            :out std_logic;
     out2019            :out std_logic;
     out2020            :out std_logic;
     out2021            :out std_logic;
     out2022            :out std_logic;
     out2023            :out std_logic;
     out2024            :out std_logic;
     out2025            :out std_logic;
     out2026            :out std_logic;
     out2027            :out std_logic;
     out2028            :out std_logic;
     out2029            :out std_logic;
     out2030            :out std_logic;
     out2031            :out std_logic;
     out2032            :out std_logic;
     out2033            :out std_logic;
     out2034            :out std_logic;
     out2035            :out std_logic;
     out2036            :out std_logic;
     out2037            :out std_logic;
     out2038            :out std_logic;
     out2039            :out std_logic;
     out2040            :out std_logic;
     out2041            :out std_logic;
     out2042            :out std_logic;
     out2043            :out std_logic;
     out2044            :out std_logic;
     out2045            :out std_logic;
     out2046            :out std_logic;
     out2047            :out std_logic;
     out2048            :out std_logic;
     out2049            :out std_logic;
     out2050            :out std_logic;
     out2051            :out std_logic;
     out2052            :out std_logic;
     out2053            :out std_logic;
     out2054            :out std_logic;
     out2055            :out std_logic;
     out2056            :out std_logic;
     out2057            :out std_logic;
     out2058            :out std_logic;
     out2059            :out std_logic;
     out2060            :out std_logic;
     out2061            :out std_logic;
     out2062            :out std_logic;
     out2063            :out std_logic;
     out2064            :out std_logic;
     out2065            :out std_logic;
     out2066            :out std_logic;
     out2067            :out std_logic;
     out2068            :out std_logic;
     out2069            :out std_logic;
     out2070            :out std_logic;
     out2071            :out std_logic;
     out2072            :out std_logic;
     out2073            :out std_logic;
     out2074            :out std_logic;
     out2075            :out std_logic;
     out2076            :out std_logic;
     out2077            :out std_logic;
     out2078            :out std_logic;
     out2079            :out std_logic;
     out2080            :out std_logic;
     out2081            :out std_logic;
     out2082            :out std_logic;
     out2083            :out std_logic;
     out2084            :out std_logic;
     out2085            :out std_logic;
     out2086            :out std_logic;
     out2087            :out std_logic;
     out2088            :out std_logic;
     out2089            :out std_logic;
     out2090            :out std_logic;
     out2091            :out std_logic;
     out2092            :out std_logic;
     out2093            :out std_logic;
     out2094            :out std_logic;
     out2095            :out std_logic;
     out2096            :out std_logic;
     out2097            :out std_logic;
     out2098            :out std_logic;
     out2099            :out std_logic;
     out2100            :out std_logic;
     out2101            :out std_logic;
     out2102            :out std_logic;
     out2103            :out std_logic;
     out2104            :out std_logic;
     out2105            :out std_logic;
     out2106            :out std_logic;
     out2107            :out std_logic;
     out2108            :out std_logic;
     out2109            :out std_logic;
     out2110            :out std_logic;
     out2111            :out std_logic;
     out2112            :out std_logic;
     out2113            :out std_logic;
     out2114            :out std_logic;
     out2115            :out std_logic;
     out2116            :out std_logic;
     out2117            :out std_logic;
     out2118            :out std_logic;
     out2119            :out std_logic;
     out2120            :out std_logic;
     out2121            :out std_logic;
     out2122            :out std_logic;
     out2123            :out std_logic;
     out2124            :out std_logic;
     out2125            :out std_logic;
     out2126            :out std_logic;
     out2127            :out std_logic;
     out2128            :out std_logic;
     out2129            :out std_logic;
     out2130            :out std_logic;
     out2131            :out std_logic;
     out2132            :out std_logic;
     out2133            :out std_logic;
     out2134            :out std_logic;
     out2135            :out std_logic;
     out2136            :out std_logic;
     out2137            :out std_logic;
     out2138            :out std_logic;
     out2139            :out std_logic;
     out2140            :out std_logic;
     out2141            :out std_logic;
     out2142            :out std_logic;
     out2143            :out std_logic;
     out2144            :out std_logic;
     out2145            :out std_logic;
     out2146            :out std_logic;
     out2147            :out std_logic;
     out2148            :out std_logic;
     out2149            :out std_logic;
     out2150            :out std_logic;
     out2151            :out std_logic;
     out2152            :out std_logic;
     out2153            :out std_logic;
     out2154            :out std_logic;
     out2155            :out std_logic;
     out2156            :out std_logic;
     out2157            :out std_logic;
     out2158            :out std_logic;
     out2159            :out std_logic;
     out2160            :out std_logic;
     out2161            :out std_logic;
     out2162            :out std_logic;
     out2163            :out std_logic;
     out2164            :out std_logic;
     out2165            :out std_logic;
     out2166            :out std_logic;
     out2167            :out std_logic;
     out2168            :out std_logic;
     out2169            :out std_logic;
     out2170            :out std_logic;
     out2171            :out std_logic;
     out2172            :out std_logic;
     out2173            :out std_logic;
     out2174            :out std_logic;
     out2175            :out std_logic;
     out2176            :out std_logic;
     out2177            :out std_logic;
     out2178            :out std_logic;
     out2179            :out std_logic;
     out2180            :out std_logic;
     out2181            :out std_logic;
     out2182            :out std_logic;
     out2183            :out std_logic;
     out2184            :out std_logic;
     out2185            :out std_logic;
     out2186            :out std_logic;
     out2187            :out std_logic;
     out2188            :out std_logic;
     out2189            :out std_logic;
     out2190            :out std_logic;
     out2191            :out std_logic;
     out2192            :out std_logic;
     out2193            :out std_logic;
     out2194            :out std_logic;
     out2195            :out std_logic;
     out2196            :out std_logic;
     out2197            :out std_logic;
     out2198            :out std_logic;
     out2199            :out std_logic;
     out2200            :out std_logic;
     out2201            :out std_logic;
     out2202            :out std_logic;
     out2203            :out std_logic;
     out2204            :out std_logic;
     out2205            :out std_logic;
     out2206            :out std_logic;
     out2207            :out std_logic;
     out2208            :out std_logic;
     out2209            :out std_logic;
     out2210            :out std_logic;
     out2211            :out std_logic;
     out2212            :out std_logic;
     out2213            :out std_logic;
     out2214            :out std_logic;
     out2215            :out std_logic;
     out2216            :out std_logic;
     out2217            :out std_logic;
     out2218            :out std_logic;
     out2219            :out std_logic;
     out2220            :out std_logic;
     out2221            :out std_logic;
     out2222            :out std_logic;
     out2223            :out std_logic;
     out2224            :out std_logic;
     out2225            :out std_logic;
     out2226            :out std_logic;
     out2227            :out std_logic;
     out2228            :out std_logic;
     out2229            :out std_logic;
     out2230            :out std_logic;
     out2231            :out std_logic;
     out2232            :out std_logic;
     out2233            :out std_logic;
     out2234            :out std_logic;
     out2235            :out std_logic;
     out2236            :out std_logic;
     out2237            :out std_logic;
     out2238            :out std_logic;
     out2239            :out std_logic;
     out2240            :out std_logic;
     out2241            :out std_logic;
     out2242            :out std_logic;
     out2243            :out std_logic;
     out2244            :out std_logic;
     out2245            :out std_logic;
     out2246            :out std_logic;
     out2247            :out std_logic;
     out2248            :out std_logic;
     out2249            :out std_logic;
     out2250            :out std_logic;
     out2251            :out std_logic;
     out2252            :out std_logic;
     out2253            :out std_logic;
     out2254            :out std_logic;
     out2255            :out std_logic;
     out2256            :out std_logic;
     out2257            :out std_logic;
     out2258            :out std_logic;
     out2259            :out std_logic;
     out2260            :out std_logic;
     out2261            :out std_logic;
     out2262            :out std_logic;
     out2263            :out std_logic;
     out2264            :out std_logic;
     out2265            :out std_logic;
     out2266            :out std_logic;
     out2267            :out std_logic;
     out2268            :out std_logic;
     out2269            :out std_logic;
     out2270            :out std_logic;
     out2271            :out std_logic;
     out2272            :out std_logic;
     out2273            :out std_logic;
     out2274            :out std_logic;
     out2275            :out std_logic;
     out2276            :out std_logic;
     out2277            :out std_logic;
     out2278            :out std_logic;
     out2279            :out std_logic;
     out2280            :out std_logic;
     out2281            :out std_logic;
     out2282            :out std_logic;
     out2283            :out std_logic;
     out2284            :out std_logic;
     out2285            :out std_logic;
     out2286            :out std_logic;
     out2287            :out std_logic;
     out2288            :out std_logic;
     out2289            :out std_logic;
     out2290            :out std_logic;
     out2291            :out std_logic;
     out2292            :out std_logic;
     out2293            :out std_logic;
     out2294            :out std_logic;
     out2295            :out std_logic;
     out2296            :out std_logic;
     out2297            :out std_logic;
     out2298            :out std_logic;
     out2299            :out std_logic;
     out2300            :out std_logic;
     out2301            :out std_logic;
     out2302            :out std_logic;
     out2303            :out std_logic;
     out2304            :out std_logic;
     end_cnt,end_vnt      :out std_logic
);
END component;

COMPONENT decision is PORT(
     clk,rst,start_pa     :in std_logic;
    iter_max      :in std_logic_vector(4 downto 0);
     x1            :in std_logic;
     x2            :in std_logic;
     x3            :in std_logic;
     x4            :in std_logic;
     x5            :in std_logic;
     x6            :in std_logic;
     x7            :in std_logic;
     x8            :in std_logic;
     x9            :in std_logic;
     x10            :in std_logic;
     x11            :in std_logic;
     x12            :in std_logic;
     x13            :in std_logic;
     x14            :in std_logic;
     x15            :in std_logic;
     x16            :in std_logic;
     x17            :in std_logic;
     x18            :in std_logic;
     x19            :in std_logic;
     x20            :in std_logic;
     x21            :in std_logic;
     x22            :in std_logic;
     x23            :in std_logic;
     x24            :in std_logic;
     x25            :in std_logic;
     x26            :in std_logic;
     x27            :in std_logic;
     x28            :in std_logic;
     x29            :in std_logic;
     x30            :in std_logic;
     x31            :in std_logic;
     x32            :in std_logic;
     x33            :in std_logic;
     x34            :in std_logic;
     x35            :in std_logic;
     x36            :in std_logic;
     x37            :in std_logic;
     x38            :in std_logic;
     x39            :in std_logic;
     x40            :in std_logic;
     x41            :in std_logic;
     x42            :in std_logic;
     x43            :in std_logic;
     x44            :in std_logic;
     x45            :in std_logic;
     x46            :in std_logic;
     x47            :in std_logic;
     x48            :in std_logic;
     x49            :in std_logic;
     x50            :in std_logic;
     x51            :in std_logic;
     x52            :in std_logic;
     x53            :in std_logic;
     x54            :in std_logic;
     x55            :in std_logic;
     x56            :in std_logic;
     x57            :in std_logic;
     x58            :in std_logic;
     x59            :in std_logic;
     x60            :in std_logic;
     x61            :in std_logic;
     x62            :in std_logic;
     x63            :in std_logic;
     x64            :in std_logic;
     x65            :in std_logic;
     x66            :in std_logic;
     x67            :in std_logic;
     x68            :in std_logic;
     x69            :in std_logic;
     x70            :in std_logic;
     x71            :in std_logic;
     x72            :in std_logic;
     x73            :in std_logic;
     x74            :in std_logic;
     x75            :in std_logic;
     x76            :in std_logic;
     x77            :in std_logic;
     x78            :in std_logic;
     x79            :in std_logic;
     x80            :in std_logic;
     x81            :in std_logic;
     x82            :in std_logic;
     x83            :in std_logic;
     x84            :in std_logic;
     x85            :in std_logic;
     x86            :in std_logic;
     x87            :in std_logic;
     x88            :in std_logic;
     x89            :in std_logic;
     x90            :in std_logic;
     x91            :in std_logic;
     x92            :in std_logic;
     x93            :in std_logic;
     x94            :in std_logic;
     x95            :in std_logic;
     x96            :in std_logic;
     x97            :in std_logic;
     x98            :in std_logic;
     x99            :in std_logic;
     x100            :in std_logic;
     x101            :in std_logic;
     x102            :in std_logic;
     x103            :in std_logic;
     x104            :in std_logic;
     x105            :in std_logic;
     x106            :in std_logic;
     x107            :in std_logic;
     x108            :in std_logic;
     x109            :in std_logic;
     x110            :in std_logic;
     x111            :in std_logic;
     x112            :in std_logic;
     x113            :in std_logic;
     x114            :in std_logic;
     x115            :in std_logic;
     x116            :in std_logic;
     x117            :in std_logic;
     x118            :in std_logic;
     x119            :in std_logic;
     x120            :in std_logic;
     x121            :in std_logic;
     x122            :in std_logic;
     x123            :in std_logic;
     x124            :in std_logic;
     x125            :in std_logic;
     x126            :in std_logic;
     x127            :in std_logic;
     x128            :in std_logic;
     x129            :in std_logic;
     x130            :in std_logic;
     x131            :in std_logic;
     x132            :in std_logic;
     x133            :in std_logic;
     x134            :in std_logic;
     x135            :in std_logic;
     x136            :in std_logic;
     x137            :in std_logic;
     x138            :in std_logic;
     x139            :in std_logic;
     x140            :in std_logic;
     x141            :in std_logic;
     x142            :in std_logic;
     x143            :in std_logic;
     x144            :in std_logic;
     x145            :in std_logic;
     x146            :in std_logic;
     x147            :in std_logic;
     x148            :in std_logic;
     x149            :in std_logic;
     x150            :in std_logic;
     x151            :in std_logic;
     x152            :in std_logic;
     x153            :in std_logic;
     x154            :in std_logic;
     x155            :in std_logic;
     x156            :in std_logic;
     x157            :in std_logic;
     x158            :in std_logic;
     x159            :in std_logic;
     x160            :in std_logic;
     x161            :in std_logic;
     x162            :in std_logic;
     x163            :in std_logic;
     x164            :in std_logic;
     x165            :in std_logic;
     x166            :in std_logic;
     x167            :in std_logic;
     x168            :in std_logic;
     x169            :in std_logic;
     x170            :in std_logic;
     x171            :in std_logic;
     x172            :in std_logic;
     x173            :in std_logic;
     x174            :in std_logic;
     x175            :in std_logic;
     x176            :in std_logic;
     x177            :in std_logic;
     x178            :in std_logic;
     x179            :in std_logic;
     x180            :in std_logic;
     x181            :in std_logic;
     x182            :in std_logic;
     x183            :in std_logic;
     x184            :in std_logic;
     x185            :in std_logic;
     x186            :in std_logic;
     x187            :in std_logic;
     x188            :in std_logic;
     x189            :in std_logic;
     x190            :in std_logic;
     x191            :in std_logic;
     x192            :in std_logic;
     x193            :in std_logic;
     x194            :in std_logic;
     x195            :in std_logic;
     x196            :in std_logic;
     x197            :in std_logic;
     x198            :in std_logic;
     x199            :in std_logic;
     x200            :in std_logic;
     x201            :in std_logic;
     x202            :in std_logic;
     x203            :in std_logic;
     x204            :in std_logic;
     x205            :in std_logic;
     x206            :in std_logic;
     x207            :in std_logic;
     x208            :in std_logic;
     x209            :in std_logic;
     x210            :in std_logic;
     x211            :in std_logic;
     x212            :in std_logic;
     x213            :in std_logic;
     x214            :in std_logic;
     x215            :in std_logic;
     x216            :in std_logic;
     x217            :in std_logic;
     x218            :in std_logic;
     x219            :in std_logic;
     x220            :in std_logic;
     x221            :in std_logic;
     x222            :in std_logic;
     x223            :in std_logic;
     x224            :in std_logic;
     x225            :in std_logic;
     x226            :in std_logic;
     x227            :in std_logic;
     x228            :in std_logic;
     x229            :in std_logic;
     x230            :in std_logic;
     x231            :in std_logic;
     x232            :in std_logic;
     x233            :in std_logic;
     x234            :in std_logic;
     x235            :in std_logic;
     x236            :in std_logic;
     x237            :in std_logic;
     x238            :in std_logic;
     x239            :in std_logic;
     x240            :in std_logic;
     x241            :in std_logic;
     x242            :in std_logic;
     x243            :in std_logic;
     x244            :in std_logic;
     x245            :in std_logic;
     x246            :in std_logic;
     x247            :in std_logic;
     x248            :in std_logic;
     x249            :in std_logic;
     x250            :in std_logic;
     x251            :in std_logic;
     x252            :in std_logic;
     x253            :in std_logic;
     x254            :in std_logic;
     x255            :in std_logic;
     x256            :in std_logic;
     x257            :in std_logic;
     x258            :in std_logic;
     x259            :in std_logic;
     x260            :in std_logic;
     x261            :in std_logic;
     x262            :in std_logic;
     x263            :in std_logic;
     x264            :in std_logic;
     x265            :in std_logic;
     x266            :in std_logic;
     x267            :in std_logic;
     x268            :in std_logic;
     x269            :in std_logic;
     x270            :in std_logic;
     x271            :in std_logic;
     x272            :in std_logic;
     x273            :in std_logic;
     x274            :in std_logic;
     x275            :in std_logic;
     x276            :in std_logic;
     x277            :in std_logic;
     x278            :in std_logic;
     x279            :in std_logic;
     x280            :in std_logic;
     x281            :in std_logic;
     x282            :in std_logic;
     x283            :in std_logic;
     x284            :in std_logic;
     x285            :in std_logic;
     x286            :in std_logic;
     x287            :in std_logic;
     x288            :in std_logic;
     x289            :in std_logic;
     x290            :in std_logic;
     x291            :in std_logic;
     x292            :in std_logic;
     x293            :in std_logic;
     x294            :in std_logic;
     x295            :in std_logic;
     x296            :in std_logic;
     x297            :in std_logic;
     x298            :in std_logic;
     x299            :in std_logic;
     x300            :in std_logic;
     x301            :in std_logic;
     x302            :in std_logic;
     x303            :in std_logic;
     x304            :in std_logic;
     x305            :in std_logic;
     x306            :in std_logic;
     x307            :in std_logic;
     x308            :in std_logic;
     x309            :in std_logic;
     x310            :in std_logic;
     x311            :in std_logic;
     x312            :in std_logic;
     x313            :in std_logic;
     x314            :in std_logic;
     x315            :in std_logic;
     x316            :in std_logic;
     x317            :in std_logic;
     x318            :in std_logic;
     x319            :in std_logic;
     x320            :in std_logic;
     x321            :in std_logic;
     x322            :in std_logic;
     x323            :in std_logic;
     x324            :in std_logic;
     x325            :in std_logic;
     x326            :in std_logic;
     x327            :in std_logic;
     x328            :in std_logic;
     x329            :in std_logic;
     x330            :in std_logic;
     x331            :in std_logic;
     x332            :in std_logic;
     x333            :in std_logic;
     x334            :in std_logic;
     x335            :in std_logic;
     x336            :in std_logic;
     x337            :in std_logic;
     x338            :in std_logic;
     x339            :in std_logic;
     x340            :in std_logic;
     x341            :in std_logic;
     x342            :in std_logic;
     x343            :in std_logic;
     x344            :in std_logic;
     x345            :in std_logic;
     x346            :in std_logic;
     x347            :in std_logic;
     x348            :in std_logic;
     x349            :in std_logic;
     x350            :in std_logic;
     x351            :in std_logic;
     x352            :in std_logic;
     x353            :in std_logic;
     x354            :in std_logic;
     x355            :in std_logic;
     x356            :in std_logic;
     x357            :in std_logic;
     x358            :in std_logic;
     x359            :in std_logic;
     x360            :in std_logic;
     x361            :in std_logic;
     x362            :in std_logic;
     x363            :in std_logic;
     x364            :in std_logic;
     x365            :in std_logic;
     x366            :in std_logic;
     x367            :in std_logic;
     x368            :in std_logic;
     x369            :in std_logic;
     x370            :in std_logic;
     x371            :in std_logic;
     x372            :in std_logic;
     x373            :in std_logic;
     x374            :in std_logic;
     x375            :in std_logic;
     x376            :in std_logic;
     x377            :in std_logic;
     x378            :in std_logic;
     x379            :in std_logic;
     x380            :in std_logic;
     x381            :in std_logic;
     x382            :in std_logic;
     x383            :in std_logic;
     x384            :in std_logic;
     x385            :in std_logic;
     x386            :in std_logic;
     x387            :in std_logic;
     x388            :in std_logic;
     x389            :in std_logic;
     x390            :in std_logic;
     x391            :in std_logic;
     x392            :in std_logic;
     x393            :in std_logic;
     x394            :in std_logic;
     x395            :in std_logic;
     x396            :in std_logic;
     x397            :in std_logic;
     x398            :in std_logic;
     x399            :in std_logic;
     x400            :in std_logic;
     x401            :in std_logic;
     x402            :in std_logic;
     x403            :in std_logic;
     x404            :in std_logic;
     x405            :in std_logic;
     x406            :in std_logic;
     x407            :in std_logic;
     x408            :in std_logic;
     x409            :in std_logic;
     x410            :in std_logic;
     x411            :in std_logic;
     x412            :in std_logic;
     x413            :in std_logic;
     x414            :in std_logic;
     x415            :in std_logic;
     x416            :in std_logic;
     x417            :in std_logic;
     x418            :in std_logic;
     x419            :in std_logic;
     x420            :in std_logic;
     x421            :in std_logic;
     x422            :in std_logic;
     x423            :in std_logic;
     x424            :in std_logic;
     x425            :in std_logic;
     x426            :in std_logic;
     x427            :in std_logic;
     x428            :in std_logic;
     x429            :in std_logic;
     x430            :in std_logic;
     x431            :in std_logic;
     x432            :in std_logic;
     x433            :in std_logic;
     x434            :in std_logic;
     x435            :in std_logic;
     x436            :in std_logic;
     x437            :in std_logic;
     x438            :in std_logic;
     x439            :in std_logic;
     x440            :in std_logic;
     x441            :in std_logic;
     x442            :in std_logic;
     x443            :in std_logic;
     x444            :in std_logic;
     x445            :in std_logic;
     x446            :in std_logic;
     x447            :in std_logic;
     x448            :in std_logic;
     x449            :in std_logic;
     x450            :in std_logic;
     x451            :in std_logic;
     x452            :in std_logic;
     x453            :in std_logic;
     x454            :in std_logic;
     x455            :in std_logic;
     x456            :in std_logic;
     x457            :in std_logic;
     x458            :in std_logic;
     x459            :in std_logic;
     x460            :in std_logic;
     x461            :in std_logic;
     x462            :in std_logic;
     x463            :in std_logic;
     x464            :in std_logic;
     x465            :in std_logic;
     x466            :in std_logic;
     x467            :in std_logic;
     x468            :in std_logic;
     x469            :in std_logic;
     x470            :in std_logic;
     x471            :in std_logic;
     x472            :in std_logic;
     x473            :in std_logic;
     x474            :in std_logic;
     x475            :in std_logic;
     x476            :in std_logic;
     x477            :in std_logic;
     x478            :in std_logic;
     x479            :in std_logic;
     x480            :in std_logic;
     x481            :in std_logic;
     x482            :in std_logic;
     x483            :in std_logic;
     x484            :in std_logic;
     x485            :in std_logic;
     x486            :in std_logic;
     x487            :in std_logic;
     x488            :in std_logic;
     x489            :in std_logic;
     x490            :in std_logic;
     x491            :in std_logic;
     x492            :in std_logic;
     x493            :in std_logic;
     x494            :in std_logic;
     x495            :in std_logic;
     x496            :in std_logic;
     x497            :in std_logic;
     x498            :in std_logic;
     x499            :in std_logic;
     x500            :in std_logic;
     x501            :in std_logic;
     x502            :in std_logic;
     x503            :in std_logic;
     x504            :in std_logic;
     x505            :in std_logic;
     x506            :in std_logic;
     x507            :in std_logic;
     x508            :in std_logic;
     x509            :in std_logic;
     x510            :in std_logic;
     x511            :in std_logic;
     x512            :in std_logic;
     x513            :in std_logic;
     x514            :in std_logic;
     x515            :in std_logic;
     x516            :in std_logic;
     x517            :in std_logic;
     x518            :in std_logic;
     x519            :in std_logic;
     x520            :in std_logic;
     x521            :in std_logic;
     x522            :in std_logic;
     x523            :in std_logic;
     x524            :in std_logic;
     x525            :in std_logic;
     x526            :in std_logic;
     x527            :in std_logic;
     x528            :in std_logic;
     x529            :in std_logic;
     x530            :in std_logic;
     x531            :in std_logic;
     x532            :in std_logic;
     x533            :in std_logic;
     x534            :in std_logic;
     x535            :in std_logic;
     x536            :in std_logic;
     x537            :in std_logic;
     x538            :in std_logic;
     x539            :in std_logic;
     x540            :in std_logic;
     x541            :in std_logic;
     x542            :in std_logic;
     x543            :in std_logic;
     x544            :in std_logic;
     x545            :in std_logic;
     x546            :in std_logic;
     x547            :in std_logic;
     x548            :in std_logic;
     x549            :in std_logic;
     x550            :in std_logic;
     x551            :in std_logic;
     x552            :in std_logic;
     x553            :in std_logic;
     x554            :in std_logic;
     x555            :in std_logic;
     x556            :in std_logic;
     x557            :in std_logic;
     x558            :in std_logic;
     x559            :in std_logic;
     x560            :in std_logic;
     x561            :in std_logic;
     x562            :in std_logic;
     x563            :in std_logic;
     x564            :in std_logic;
     x565            :in std_logic;
     x566            :in std_logic;
     x567            :in std_logic;
     x568            :in std_logic;
     x569            :in std_logic;
     x570            :in std_logic;
     x571            :in std_logic;
     x572            :in std_logic;
     x573            :in std_logic;
     x574            :in std_logic;
     x575            :in std_logic;
     x576            :in std_logic;
     x577            :in std_logic;
     x578            :in std_logic;
     x579            :in std_logic;
     x580            :in std_logic;
     x581            :in std_logic;
     x582            :in std_logic;
     x583            :in std_logic;
     x584            :in std_logic;
     x585            :in std_logic;
     x586            :in std_logic;
     x587            :in std_logic;
     x588            :in std_logic;
     x589            :in std_logic;
     x590            :in std_logic;
     x591            :in std_logic;
     x592            :in std_logic;
     x593            :in std_logic;
     x594            :in std_logic;
     x595            :in std_logic;
     x596            :in std_logic;
     x597            :in std_logic;
     x598            :in std_logic;
     x599            :in std_logic;
     x600            :in std_logic;
     x601            :in std_logic;
     x602            :in std_logic;
     x603            :in std_logic;
     x604            :in std_logic;
     x605            :in std_logic;
     x606            :in std_logic;
     x607            :in std_logic;
     x608            :in std_logic;
     x609            :in std_logic;
     x610            :in std_logic;
     x611            :in std_logic;
     x612            :in std_logic;
     x613            :in std_logic;
     x614            :in std_logic;
     x615            :in std_logic;
     x616            :in std_logic;
     x617            :in std_logic;
     x618            :in std_logic;
     x619            :in std_logic;
     x620            :in std_logic;
     x621            :in std_logic;
     x622            :in std_logic;
     x623            :in std_logic;
     x624            :in std_logic;
     x625            :in std_logic;
     x626            :in std_logic;
     x627            :in std_logic;
     x628            :in std_logic;
     x629            :in std_logic;
     x630            :in std_logic;
     x631            :in std_logic;
     x632            :in std_logic;
     x633            :in std_logic;
     x634            :in std_logic;
     x635            :in std_logic;
     x636            :in std_logic;
     x637            :in std_logic;
     x638            :in std_logic;
     x639            :in std_logic;
     x640            :in std_logic;
     x641            :in std_logic;
     x642            :in std_logic;
     x643            :in std_logic;
     x644            :in std_logic;
     x645            :in std_logic;
     x646            :in std_logic;
     x647            :in std_logic;
     x648            :in std_logic;
     x649            :in std_logic;
     x650            :in std_logic;
     x651            :in std_logic;
     x652            :in std_logic;
     x653            :in std_logic;
     x654            :in std_logic;
     x655            :in std_logic;
     x656            :in std_logic;
     x657            :in std_logic;
     x658            :in std_logic;
     x659            :in std_logic;
     x660            :in std_logic;
     x661            :in std_logic;
     x662            :in std_logic;
     x663            :in std_logic;
     x664            :in std_logic;
     x665            :in std_logic;
     x666            :in std_logic;
     x667            :in std_logic;
     x668            :in std_logic;
     x669            :in std_logic;
     x670            :in std_logic;
     x671            :in std_logic;
     x672            :in std_logic;
     x673            :in std_logic;
     x674            :in std_logic;
     x675            :in std_logic;
     x676            :in std_logic;
     x677            :in std_logic;
     x678            :in std_logic;
     x679            :in std_logic;
     x680            :in std_logic;
     x681            :in std_logic;
     x682            :in std_logic;
     x683            :in std_logic;
     x684            :in std_logic;
     x685            :in std_logic;
     x686            :in std_logic;
     x687            :in std_logic;
     x688            :in std_logic;
     x689            :in std_logic;
     x690            :in std_logic;
     x691            :in std_logic;
     x692            :in std_logic;
     x693            :in std_logic;
     x694            :in std_logic;
     x695            :in std_logic;
     x696            :in std_logic;
     x697            :in std_logic;
     x698            :in std_logic;
     x699            :in std_logic;
     x700            :in std_logic;
     x701            :in std_logic;
     x702            :in std_logic;
     x703            :in std_logic;
     x704            :in std_logic;
     x705            :in std_logic;
     x706            :in std_logic;
     x707            :in std_logic;
     x708            :in std_logic;
     x709            :in std_logic;
     x710            :in std_logic;
     x711            :in std_logic;
     x712            :in std_logic;
     x713            :in std_logic;
     x714            :in std_logic;
     x715            :in std_logic;
     x716            :in std_logic;
     x717            :in std_logic;
     x718            :in std_logic;
     x719            :in std_logic;
     x720            :in std_logic;
     x721            :in std_logic;
     x722            :in std_logic;
     x723            :in std_logic;
     x724            :in std_logic;
     x725            :in std_logic;
     x726            :in std_logic;
     x727            :in std_logic;
     x728            :in std_logic;
     x729            :in std_logic;
     x730            :in std_logic;
     x731            :in std_logic;
     x732            :in std_logic;
     x733            :in std_logic;
     x734            :in std_logic;
     x735            :in std_logic;
     x736            :in std_logic;
     x737            :in std_logic;
     x738            :in std_logic;
     x739            :in std_logic;
     x740            :in std_logic;
     x741            :in std_logic;
     x742            :in std_logic;
     x743            :in std_logic;
     x744            :in std_logic;
     x745            :in std_logic;
     x746            :in std_logic;
     x747            :in std_logic;
     x748            :in std_logic;
     x749            :in std_logic;
     x750            :in std_logic;
     x751            :in std_logic;
     x752            :in std_logic;
     x753            :in std_logic;
     x754            :in std_logic;
     x755            :in std_logic;
     x756            :in std_logic;
     x757            :in std_logic;
     x758            :in std_logic;
     x759            :in std_logic;
     x760            :in std_logic;
     x761            :in std_logic;
     x762            :in std_logic;
     x763            :in std_logic;
     x764            :in std_logic;
     x765            :in std_logic;
     x766            :in std_logic;
     x767            :in std_logic;
     x768            :in std_logic;
     x769            :in std_logic;
     x770            :in std_logic;
     x771            :in std_logic;
     x772            :in std_logic;
     x773            :in std_logic;
     x774            :in std_logic;
     x775            :in std_logic;
     x776            :in std_logic;
     x777            :in std_logic;
     x778            :in std_logic;
     x779            :in std_logic;
     x780            :in std_logic;
     x781            :in std_logic;
     x782            :in std_logic;
     x783            :in std_logic;
     x784            :in std_logic;
     x785            :in std_logic;
     x786            :in std_logic;
     x787            :in std_logic;
     x788            :in std_logic;
     x789            :in std_logic;
     x790            :in std_logic;
     x791            :in std_logic;
     x792            :in std_logic;
     x793            :in std_logic;
     x794            :in std_logic;
     x795            :in std_logic;
     x796            :in std_logic;
     x797            :in std_logic;
     x798            :in std_logic;
     x799            :in std_logic;
     x800            :in std_logic;
     x801            :in std_logic;
     x802            :in std_logic;
     x803            :in std_logic;
     x804            :in std_logic;
     x805            :in std_logic;
     x806            :in std_logic;
     x807            :in std_logic;
     x808            :in std_logic;
     x809            :in std_logic;
     x810            :in std_logic;
     x811            :in std_logic;
     x812            :in std_logic;
     x813            :in std_logic;
     x814            :in std_logic;
     x815            :in std_logic;
     x816            :in std_logic;
     x817            :in std_logic;
     x818            :in std_logic;
     x819            :in std_logic;
     x820            :in std_logic;
     x821            :in std_logic;
     x822            :in std_logic;
     x823            :in std_logic;
     x824            :in std_logic;
     x825            :in std_logic;
     x826            :in std_logic;
     x827            :in std_logic;
     x828            :in std_logic;
     x829            :in std_logic;
     x830            :in std_logic;
     x831            :in std_logic;
     x832            :in std_logic;
     x833            :in std_logic;
     x834            :in std_logic;
     x835            :in std_logic;
     x836            :in std_logic;
     x837            :in std_logic;
     x838            :in std_logic;
     x839            :in std_logic;
     x840            :in std_logic;
     x841            :in std_logic;
     x842            :in std_logic;
     x843            :in std_logic;
     x844            :in std_logic;
     x845            :in std_logic;
     x846            :in std_logic;
     x847            :in std_logic;
     x848            :in std_logic;
     x849            :in std_logic;
     x850            :in std_logic;
     x851            :in std_logic;
     x852            :in std_logic;
     x853            :in std_logic;
     x854            :in std_logic;
     x855            :in std_logic;
     x856            :in std_logic;
     x857            :in std_logic;
     x858            :in std_logic;
     x859            :in std_logic;
     x860            :in std_logic;
     x861            :in std_logic;
     x862            :in std_logic;
     x863            :in std_logic;
     x864            :in std_logic;
     x865            :in std_logic;
     x866            :in std_logic;
     x867            :in std_logic;
     x868            :in std_logic;
     x869            :in std_logic;
     x870            :in std_logic;
     x871            :in std_logic;
     x872            :in std_logic;
     x873            :in std_logic;
     x874            :in std_logic;
     x875            :in std_logic;
     x876            :in std_logic;
     x877            :in std_logic;
     x878            :in std_logic;
     x879            :in std_logic;
     x880            :in std_logic;
     x881            :in std_logic;
     x882            :in std_logic;
     x883            :in std_logic;
     x884            :in std_logic;
     x885            :in std_logic;
     x886            :in std_logic;
     x887            :in std_logic;
     x888            :in std_logic;
     x889            :in std_logic;
     x890            :in std_logic;
     x891            :in std_logic;
     x892            :in std_logic;
     x893            :in std_logic;
     x894            :in std_logic;
     x895            :in std_logic;
     x896            :in std_logic;
     x897            :in std_logic;
     x898            :in std_logic;
     x899            :in std_logic;
     x900            :in std_logic;
     x901            :in std_logic;
     x902            :in std_logic;
     x903            :in std_logic;
     x904            :in std_logic;
     x905            :in std_logic;
     x906            :in std_logic;
     x907            :in std_logic;
     x908            :in std_logic;
     x909            :in std_logic;
     x910            :in std_logic;
     x911            :in std_logic;
     x912            :in std_logic;
     x913            :in std_logic;
     x914            :in std_logic;
     x915            :in std_logic;
     x916            :in std_logic;
     x917            :in std_logic;
     x918            :in std_logic;
     x919            :in std_logic;
     x920            :in std_logic;
     x921            :in std_logic;
     x922            :in std_logic;
     x923            :in std_logic;
     x924            :in std_logic;
     x925            :in std_logic;
     x926            :in std_logic;
     x927            :in std_logic;
     x928            :in std_logic;
     x929            :in std_logic;
     x930            :in std_logic;
     x931            :in std_logic;
     x932            :in std_logic;
     x933            :in std_logic;
     x934            :in std_logic;
     x935            :in std_logic;
     x936            :in std_logic;
     x937            :in std_logic;
     x938            :in std_logic;
     x939            :in std_logic;
     x940            :in std_logic;
     x941            :in std_logic;
     x942            :in std_logic;
     x943            :in std_logic;
     x944            :in std_logic;
     x945            :in std_logic;
     x946            :in std_logic;
     x947            :in std_logic;
     x948            :in std_logic;
     x949            :in std_logic;
     x950            :in std_logic;
     x951            :in std_logic;
     x952            :in std_logic;
     x953            :in std_logic;
     x954            :in std_logic;
     x955            :in std_logic;
     x956            :in std_logic;
     x957            :in std_logic;
     x958            :in std_logic;
     x959            :in std_logic;
     x960            :in std_logic;
     x961            :in std_logic;
     x962            :in std_logic;
     x963            :in std_logic;
     x964            :in std_logic;
     x965            :in std_logic;
     x966            :in std_logic;
     x967            :in std_logic;
     x968            :in std_logic;
     x969            :in std_logic;
     x970            :in std_logic;
     x971            :in std_logic;
     x972            :in std_logic;
     x973            :in std_logic;
     x974            :in std_logic;
     x975            :in std_logic;
     x976            :in std_logic;
     x977            :in std_logic;
     x978            :in std_logic;
     x979            :in std_logic;
     x980            :in std_logic;
     x981            :in std_logic;
     x982            :in std_logic;
     x983            :in std_logic;
     x984            :in std_logic;
     x985            :in std_logic;
     x986            :in std_logic;
     x987            :in std_logic;
     x988            :in std_logic;
     x989            :in std_logic;
     x990            :in std_logic;
     x991            :in std_logic;
     x992            :in std_logic;
     x993            :in std_logic;
     x994            :in std_logic;
     x995            :in std_logic;
     x996            :in std_logic;
     x997            :in std_logic;
     x998            :in std_logic;
     x999            :in std_logic;
     x1000            :in std_logic;
     x1001            :in std_logic;
     x1002            :in std_logic;
     x1003            :in std_logic;
     x1004            :in std_logic;
     x1005            :in std_logic;
     x1006            :in std_logic;
     x1007            :in std_logic;
     x1008            :in std_logic;
     x1009            :in std_logic;
     x1010            :in std_logic;
     x1011            :in std_logic;
     x1012            :in std_logic;
     x1013            :in std_logic;
     x1014            :in std_logic;
     x1015            :in std_logic;
     x1016            :in std_logic;
     x1017            :in std_logic;
     x1018            :in std_logic;
     x1019            :in std_logic;
     x1020            :in std_logic;
     x1021            :in std_logic;
     x1022            :in std_logic;
     x1023            :in std_logic;
     x1024            :in std_logic;
     x1025            :in std_logic;
     x1026            :in std_logic;
     x1027            :in std_logic;
     x1028            :in std_logic;
     x1029            :in std_logic;
     x1030            :in std_logic;
     x1031            :in std_logic;
     x1032            :in std_logic;
     x1033            :in std_logic;
     x1034            :in std_logic;
     x1035            :in std_logic;
     x1036            :in std_logic;
     x1037            :in std_logic;
     x1038            :in std_logic;
     x1039            :in std_logic;
     x1040            :in std_logic;
     x1041            :in std_logic;
     x1042            :in std_logic;
     x1043            :in std_logic;
     x1044            :in std_logic;
     x1045            :in std_logic;
     x1046            :in std_logic;
     x1047            :in std_logic;
     x1048            :in std_logic;
     x1049            :in std_logic;
     x1050            :in std_logic;
     x1051            :in std_logic;
     x1052            :in std_logic;
     x1053            :in std_logic;
     x1054            :in std_logic;
     x1055            :in std_logic;
     x1056            :in std_logic;
     x1057            :in std_logic;
     x1058            :in std_logic;
     x1059            :in std_logic;
     x1060            :in std_logic;
     x1061            :in std_logic;
     x1062            :in std_logic;
     x1063            :in std_logic;
     x1064            :in std_logic;
     x1065            :in std_logic;
     x1066            :in std_logic;
     x1067            :in std_logic;
     x1068            :in std_logic;
     x1069            :in std_logic;
     x1070            :in std_logic;
     x1071            :in std_logic;
     x1072            :in std_logic;
     x1073            :in std_logic;
     x1074            :in std_logic;
     x1075            :in std_logic;
     x1076            :in std_logic;
     x1077            :in std_logic;
     x1078            :in std_logic;
     x1079            :in std_logic;
     x1080            :in std_logic;
     x1081            :in std_logic;
     x1082            :in std_logic;
     x1083            :in std_logic;
     x1084            :in std_logic;
     x1085            :in std_logic;
     x1086            :in std_logic;
     x1087            :in std_logic;
     x1088            :in std_logic;
     x1089            :in std_logic;
     x1090            :in std_logic;
     x1091            :in std_logic;
     x1092            :in std_logic;
     x1093            :in std_logic;
     x1094            :in std_logic;
     x1095            :in std_logic;
     x1096            :in std_logic;
     x1097            :in std_logic;
     x1098            :in std_logic;
     x1099            :in std_logic;
     x1100            :in std_logic;
     x1101            :in std_logic;
     x1102            :in std_logic;
     x1103            :in std_logic;
     x1104            :in std_logic;
     x1105            :in std_logic;
     x1106            :in std_logic;
     x1107            :in std_logic;
     x1108            :in std_logic;
     x1109            :in std_logic;
     x1110            :in std_logic;
     x1111            :in std_logic;
     x1112            :in std_logic;
     x1113            :in std_logic;
     x1114            :in std_logic;
     x1115            :in std_logic;
     x1116            :in std_logic;
     x1117            :in std_logic;
     x1118            :in std_logic;
     x1119            :in std_logic;
     x1120            :in std_logic;
     x1121            :in std_logic;
     x1122            :in std_logic;
     x1123            :in std_logic;
     x1124            :in std_logic;
     x1125            :in std_logic;
     x1126            :in std_logic;
     x1127            :in std_logic;
     x1128            :in std_logic;
     x1129            :in std_logic;
     x1130            :in std_logic;
     x1131            :in std_logic;
     x1132            :in std_logic;
     x1133            :in std_logic;
     x1134            :in std_logic;
     x1135            :in std_logic;
     x1136            :in std_logic;
     x1137            :in std_logic;
     x1138            :in std_logic;
     x1139            :in std_logic;
     x1140            :in std_logic;
     x1141            :in std_logic;
     x1142            :in std_logic;
     x1143            :in std_logic;
     x1144            :in std_logic;
     x1145            :in std_logic;
     x1146            :in std_logic;
     x1147            :in std_logic;
     x1148            :in std_logic;
     x1149            :in std_logic;
     x1150            :in std_logic;
     x1151            :in std_logic;
     x1152            :in std_logic;
     x1153            :in std_logic;
     x1154            :in std_logic;
     x1155            :in std_logic;
     x1156            :in std_logic;
     x1157            :in std_logic;
     x1158            :in std_logic;
     x1159            :in std_logic;
     x1160            :in std_logic;
     x1161            :in std_logic;
     x1162            :in std_logic;
     x1163            :in std_logic;
     x1164            :in std_logic;
     x1165            :in std_logic;
     x1166            :in std_logic;
     x1167            :in std_logic;
     x1168            :in std_logic;
     x1169            :in std_logic;
     x1170            :in std_logic;
     x1171            :in std_logic;
     x1172            :in std_logic;
     x1173            :in std_logic;
     x1174            :in std_logic;
     x1175            :in std_logic;
     x1176            :in std_logic;
     x1177            :in std_logic;
     x1178            :in std_logic;
     x1179            :in std_logic;
     x1180            :in std_logic;
     x1181            :in std_logic;
     x1182            :in std_logic;
     x1183            :in std_logic;
     x1184            :in std_logic;
     x1185            :in std_logic;
     x1186            :in std_logic;
     x1187            :in std_logic;
     x1188            :in std_logic;
     x1189            :in std_logic;
     x1190            :in std_logic;
     x1191            :in std_logic;
     x1192            :in std_logic;
     x1193            :in std_logic;
     x1194            :in std_logic;
     x1195            :in std_logic;
     x1196            :in std_logic;
     x1197            :in std_logic;
     x1198            :in std_logic;
     x1199            :in std_logic;
     x1200            :in std_logic;
     x1201            :in std_logic;
     x1202            :in std_logic;
     x1203            :in std_logic;
     x1204            :in std_logic;
     x1205            :in std_logic;
     x1206            :in std_logic;
     x1207            :in std_logic;
     x1208            :in std_logic;
     x1209            :in std_logic;
     x1210            :in std_logic;
     x1211            :in std_logic;
     x1212            :in std_logic;
     x1213            :in std_logic;
     x1214            :in std_logic;
     x1215            :in std_logic;
     x1216            :in std_logic;
     x1217            :in std_logic;
     x1218            :in std_logic;
     x1219            :in std_logic;
     x1220            :in std_logic;
     x1221            :in std_logic;
     x1222            :in std_logic;
     x1223            :in std_logic;
     x1224            :in std_logic;
     x1225            :in std_logic;
     x1226            :in std_logic;
     x1227            :in std_logic;
     x1228            :in std_logic;
     x1229            :in std_logic;
     x1230            :in std_logic;
     x1231            :in std_logic;
     x1232            :in std_logic;
     x1233            :in std_logic;
     x1234            :in std_logic;
     x1235            :in std_logic;
     x1236            :in std_logic;
     x1237            :in std_logic;
     x1238            :in std_logic;
     x1239            :in std_logic;
     x1240            :in std_logic;
     x1241            :in std_logic;
     x1242            :in std_logic;
     x1243            :in std_logic;
     x1244            :in std_logic;
     x1245            :in std_logic;
     x1246            :in std_logic;
     x1247            :in std_logic;
     x1248            :in std_logic;
     x1249            :in std_logic;
     x1250            :in std_logic;
     x1251            :in std_logic;
     x1252            :in std_logic;
     x1253            :in std_logic;
     x1254            :in std_logic;
     x1255            :in std_logic;
     x1256            :in std_logic;
     x1257            :in std_logic;
     x1258            :in std_logic;
     x1259            :in std_logic;
     x1260            :in std_logic;
     x1261            :in std_logic;
     x1262            :in std_logic;
     x1263            :in std_logic;
     x1264            :in std_logic;
     x1265            :in std_logic;
     x1266            :in std_logic;
     x1267            :in std_logic;
     x1268            :in std_logic;
     x1269            :in std_logic;
     x1270            :in std_logic;
     x1271            :in std_logic;
     x1272            :in std_logic;
     x1273            :in std_logic;
     x1274            :in std_logic;
     x1275            :in std_logic;
     x1276            :in std_logic;
     x1277            :in std_logic;
     x1278            :in std_logic;
     x1279            :in std_logic;
     x1280            :in std_logic;
     x1281            :in std_logic;
     x1282            :in std_logic;
     x1283            :in std_logic;
     x1284            :in std_logic;
     x1285            :in std_logic;
     x1286            :in std_logic;
     x1287            :in std_logic;
     x1288            :in std_logic;
     x1289            :in std_logic;
     x1290            :in std_logic;
     x1291            :in std_logic;
     x1292            :in std_logic;
     x1293            :in std_logic;
     x1294            :in std_logic;
     x1295            :in std_logic;
     x1296            :in std_logic;
     x1297            :in std_logic;
     x1298            :in std_logic;
     x1299            :in std_logic;
     x1300            :in std_logic;
     x1301            :in std_logic;
     x1302            :in std_logic;
     x1303            :in std_logic;
     x1304            :in std_logic;
     x1305            :in std_logic;
     x1306            :in std_logic;
     x1307            :in std_logic;
     x1308            :in std_logic;
     x1309            :in std_logic;
     x1310            :in std_logic;
     x1311            :in std_logic;
     x1312            :in std_logic;
     x1313            :in std_logic;
     x1314            :in std_logic;
     x1315            :in std_logic;
     x1316            :in std_logic;
     x1317            :in std_logic;
     x1318            :in std_logic;
     x1319            :in std_logic;
     x1320            :in std_logic;
     x1321            :in std_logic;
     x1322            :in std_logic;
     x1323            :in std_logic;
     x1324            :in std_logic;
     x1325            :in std_logic;
     x1326            :in std_logic;
     x1327            :in std_logic;
     x1328            :in std_logic;
     x1329            :in std_logic;
     x1330            :in std_logic;
     x1331            :in std_logic;
     x1332            :in std_logic;
     x1333            :in std_logic;
     x1334            :in std_logic;
     x1335            :in std_logic;
     x1336            :in std_logic;
     x1337            :in std_logic;
     x1338            :in std_logic;
     x1339            :in std_logic;
     x1340            :in std_logic;
     x1341            :in std_logic;
     x1342            :in std_logic;
     x1343            :in std_logic;
     x1344            :in std_logic;
     x1345            :in std_logic;
     x1346            :in std_logic;
     x1347            :in std_logic;
     x1348            :in std_logic;
     x1349            :in std_logic;
     x1350            :in std_logic;
     x1351            :in std_logic;
     x1352            :in std_logic;
     x1353            :in std_logic;
     x1354            :in std_logic;
     x1355            :in std_logic;
     x1356            :in std_logic;
     x1357            :in std_logic;
     x1358            :in std_logic;
     x1359            :in std_logic;
     x1360            :in std_logic;
     x1361            :in std_logic;
     x1362            :in std_logic;
     x1363            :in std_logic;
     x1364            :in std_logic;
     x1365            :in std_logic;
     x1366            :in std_logic;
     x1367            :in std_logic;
     x1368            :in std_logic;
     x1369            :in std_logic;
     x1370            :in std_logic;
     x1371            :in std_logic;
     x1372            :in std_logic;
     x1373            :in std_logic;
     x1374            :in std_logic;
     x1375            :in std_logic;
     x1376            :in std_logic;
     x1377            :in std_logic;
     x1378            :in std_logic;
     x1379            :in std_logic;
     x1380            :in std_logic;
     x1381            :in std_logic;
     x1382            :in std_logic;
     x1383            :in std_logic;
     x1384            :in std_logic;
     x1385            :in std_logic;
     x1386            :in std_logic;
     x1387            :in std_logic;
     x1388            :in std_logic;
     x1389            :in std_logic;
     x1390            :in std_logic;
     x1391            :in std_logic;
     x1392            :in std_logic;
     x1393            :in std_logic;
     x1394            :in std_logic;
     x1395            :in std_logic;
     x1396            :in std_logic;
     x1397            :in std_logic;
     x1398            :in std_logic;
     x1399            :in std_logic;
     x1400            :in std_logic;
     x1401            :in std_logic;
     x1402            :in std_logic;
     x1403            :in std_logic;
     x1404            :in std_logic;
     x1405            :in std_logic;
     x1406            :in std_logic;
     x1407            :in std_logic;
     x1408            :in std_logic;
     x1409            :in std_logic;
     x1410            :in std_logic;
     x1411            :in std_logic;
     x1412            :in std_logic;
     x1413            :in std_logic;
     x1414            :in std_logic;
     x1415            :in std_logic;
     x1416            :in std_logic;
     x1417            :in std_logic;
     x1418            :in std_logic;
     x1419            :in std_logic;
     x1420            :in std_logic;
     x1421            :in std_logic;
     x1422            :in std_logic;
     x1423            :in std_logic;
     x1424            :in std_logic;
     x1425            :in std_logic;
     x1426            :in std_logic;
     x1427            :in std_logic;
     x1428            :in std_logic;
     x1429            :in std_logic;
     x1430            :in std_logic;
     x1431            :in std_logic;
     x1432            :in std_logic;
     x1433            :in std_logic;
     x1434            :in std_logic;
     x1435            :in std_logic;
     x1436            :in std_logic;
     x1437            :in std_logic;
     x1438            :in std_logic;
     x1439            :in std_logic;
     x1440            :in std_logic;
     x1441            :in std_logic;
     x1442            :in std_logic;
     x1443            :in std_logic;
     x1444            :in std_logic;
     x1445            :in std_logic;
     x1446            :in std_logic;
     x1447            :in std_logic;
     x1448            :in std_logic;
     x1449            :in std_logic;
     x1450            :in std_logic;
     x1451            :in std_logic;
     x1452            :in std_logic;
     x1453            :in std_logic;
     x1454            :in std_logic;
     x1455            :in std_logic;
     x1456            :in std_logic;
     x1457            :in std_logic;
     x1458            :in std_logic;
     x1459            :in std_logic;
     x1460            :in std_logic;
     x1461            :in std_logic;
     x1462            :in std_logic;
     x1463            :in std_logic;
     x1464            :in std_logic;
     x1465            :in std_logic;
     x1466            :in std_logic;
     x1467            :in std_logic;
     x1468            :in std_logic;
     x1469            :in std_logic;
     x1470            :in std_logic;
     x1471            :in std_logic;
     x1472            :in std_logic;
     x1473            :in std_logic;
     x1474            :in std_logic;
     x1475            :in std_logic;
     x1476            :in std_logic;
     x1477            :in std_logic;
     x1478            :in std_logic;
     x1479            :in std_logic;
     x1480            :in std_logic;
     x1481            :in std_logic;
     x1482            :in std_logic;
     x1483            :in std_logic;
     x1484            :in std_logic;
     x1485            :in std_logic;
     x1486            :in std_logic;
     x1487            :in std_logic;
     x1488            :in std_logic;
     x1489            :in std_logic;
     x1490            :in std_logic;
     x1491            :in std_logic;
     x1492            :in std_logic;
     x1493            :in std_logic;
     x1494            :in std_logic;
     x1495            :in std_logic;
     x1496            :in std_logic;
     x1497            :in std_logic;
     x1498            :in std_logic;
     x1499            :in std_logic;
     x1500            :in std_logic;
     x1501            :in std_logic;
     x1502            :in std_logic;
     x1503            :in std_logic;
     x1504            :in std_logic;
     x1505            :in std_logic;
     x1506            :in std_logic;
     x1507            :in std_logic;
     x1508            :in std_logic;
     x1509            :in std_logic;
     x1510            :in std_logic;
     x1511            :in std_logic;
     x1512            :in std_logic;
     x1513            :in std_logic;
     x1514            :in std_logic;
     x1515            :in std_logic;
     x1516            :in std_logic;
     x1517            :in std_logic;
     x1518            :in std_logic;
     x1519            :in std_logic;
     x1520            :in std_logic;
     x1521            :in std_logic;
     x1522            :in std_logic;
     x1523            :in std_logic;
     x1524            :in std_logic;
     x1525            :in std_logic;
     x1526            :in std_logic;
     x1527            :in std_logic;
     x1528            :in std_logic;
     x1529            :in std_logic;
     x1530            :in std_logic;
     x1531            :in std_logic;
     x1532            :in std_logic;
     x1533            :in std_logic;
     x1534            :in std_logic;
     x1535            :in std_logic;
     x1536            :in std_logic;
     x1537            :in std_logic;
     x1538            :in std_logic;
     x1539            :in std_logic;
     x1540            :in std_logic;
     x1541            :in std_logic;
     x1542            :in std_logic;
     x1543            :in std_logic;
     x1544            :in std_logic;
     x1545            :in std_logic;
     x1546            :in std_logic;
     x1547            :in std_logic;
     x1548            :in std_logic;
     x1549            :in std_logic;
     x1550            :in std_logic;
     x1551            :in std_logic;
     x1552            :in std_logic;
     x1553            :in std_logic;
     x1554            :in std_logic;
     x1555            :in std_logic;
     x1556            :in std_logic;
     x1557            :in std_logic;
     x1558            :in std_logic;
     x1559            :in std_logic;
     x1560            :in std_logic;
     x1561            :in std_logic;
     x1562            :in std_logic;
     x1563            :in std_logic;
     x1564            :in std_logic;
     x1565            :in std_logic;
     x1566            :in std_logic;
     x1567            :in std_logic;
     x1568            :in std_logic;
     x1569            :in std_logic;
     x1570            :in std_logic;
     x1571            :in std_logic;
     x1572            :in std_logic;
     x1573            :in std_logic;
     x1574            :in std_logic;
     x1575            :in std_logic;
     x1576            :in std_logic;
     x1577            :in std_logic;
     x1578            :in std_logic;
     x1579            :in std_logic;
     x1580            :in std_logic;
     x1581            :in std_logic;
     x1582            :in std_logic;
     x1583            :in std_logic;
     x1584            :in std_logic;
     x1585            :in std_logic;
     x1586            :in std_logic;
     x1587            :in std_logic;
     x1588            :in std_logic;
     x1589            :in std_logic;
     x1590            :in std_logic;
     x1591            :in std_logic;
     x1592            :in std_logic;
     x1593            :in std_logic;
     x1594            :in std_logic;
     x1595            :in std_logic;
     x1596            :in std_logic;
     x1597            :in std_logic;
     x1598            :in std_logic;
     x1599            :in std_logic;
     x1600            :in std_logic;
     x1601            :in std_logic;
     x1602            :in std_logic;
     x1603            :in std_logic;
     x1604            :in std_logic;
     x1605            :in std_logic;
     x1606            :in std_logic;
     x1607            :in std_logic;
     x1608            :in std_logic;
     x1609            :in std_logic;
     x1610            :in std_logic;
     x1611            :in std_logic;
     x1612            :in std_logic;
     x1613            :in std_logic;
     x1614            :in std_logic;
     x1615            :in std_logic;
     x1616            :in std_logic;
     x1617            :in std_logic;
     x1618            :in std_logic;
     x1619            :in std_logic;
     x1620            :in std_logic;
     x1621            :in std_logic;
     x1622            :in std_logic;
     x1623            :in std_logic;
     x1624            :in std_logic;
     x1625            :in std_logic;
     x1626            :in std_logic;
     x1627            :in std_logic;
     x1628            :in std_logic;
     x1629            :in std_logic;
     x1630            :in std_logic;
     x1631            :in std_logic;
     x1632            :in std_logic;
     x1633            :in std_logic;
     x1634            :in std_logic;
     x1635            :in std_logic;
     x1636            :in std_logic;
     x1637            :in std_logic;
     x1638            :in std_logic;
     x1639            :in std_logic;
     x1640            :in std_logic;
     x1641            :in std_logic;
     x1642            :in std_logic;
     x1643            :in std_logic;
     x1644            :in std_logic;
     x1645            :in std_logic;
     x1646            :in std_logic;
     x1647            :in std_logic;
     x1648            :in std_logic;
     x1649            :in std_logic;
     x1650            :in std_logic;
     x1651            :in std_logic;
     x1652            :in std_logic;
     x1653            :in std_logic;
     x1654            :in std_logic;
     x1655            :in std_logic;
     x1656            :in std_logic;
     x1657            :in std_logic;
     x1658            :in std_logic;
     x1659            :in std_logic;
     x1660            :in std_logic;
     x1661            :in std_logic;
     x1662            :in std_logic;
     x1663            :in std_logic;
     x1664            :in std_logic;
     x1665            :in std_logic;
     x1666            :in std_logic;
     x1667            :in std_logic;
     x1668            :in std_logic;
     x1669            :in std_logic;
     x1670            :in std_logic;
     x1671            :in std_logic;
     x1672            :in std_logic;
     x1673            :in std_logic;
     x1674            :in std_logic;
     x1675            :in std_logic;
     x1676            :in std_logic;
     x1677            :in std_logic;
     x1678            :in std_logic;
     x1679            :in std_logic;
     x1680            :in std_logic;
     x1681            :in std_logic;
     x1682            :in std_logic;
     x1683            :in std_logic;
     x1684            :in std_logic;
     x1685            :in std_logic;
     x1686            :in std_logic;
     x1687            :in std_logic;
     x1688            :in std_logic;
     x1689            :in std_logic;
     x1690            :in std_logic;
     x1691            :in std_logic;
     x1692            :in std_logic;
     x1693            :in std_logic;
     x1694            :in std_logic;
     x1695            :in std_logic;
     x1696            :in std_logic;
     x1697            :in std_logic;
     x1698            :in std_logic;
     x1699            :in std_logic;
     x1700            :in std_logic;
     x1701            :in std_logic;
     x1702            :in std_logic;
     x1703            :in std_logic;
     x1704            :in std_logic;
     x1705            :in std_logic;
     x1706            :in std_logic;
     x1707            :in std_logic;
     x1708            :in std_logic;
     x1709            :in std_logic;
     x1710            :in std_logic;
     x1711            :in std_logic;
     x1712            :in std_logic;
     x1713            :in std_logic;
     x1714            :in std_logic;
     x1715            :in std_logic;
     x1716            :in std_logic;
     x1717            :in std_logic;
     x1718            :in std_logic;
     x1719            :in std_logic;
     x1720            :in std_logic;
     x1721            :in std_logic;
     x1722            :in std_logic;
     x1723            :in std_logic;
     x1724            :in std_logic;
     x1725            :in std_logic;
     x1726            :in std_logic;
     x1727            :in std_logic;
     x1728            :in std_logic;
     x1729            :in std_logic;
     x1730            :in std_logic;
     x1731            :in std_logic;
     x1732            :in std_logic;
     x1733            :in std_logic;
     x1734            :in std_logic;
     x1735            :in std_logic;
     x1736            :in std_logic;
     x1737            :in std_logic;
     x1738            :in std_logic;
     x1739            :in std_logic;
     x1740            :in std_logic;
     x1741            :in std_logic;
     x1742            :in std_logic;
     x1743            :in std_logic;
     x1744            :in std_logic;
     x1745            :in std_logic;
     x1746            :in std_logic;
     x1747            :in std_logic;
     x1748            :in std_logic;
     x1749            :in std_logic;
     x1750            :in std_logic;
     x1751            :in std_logic;
     x1752            :in std_logic;
     x1753            :in std_logic;
     x1754            :in std_logic;
     x1755            :in std_logic;
     x1756            :in std_logic;
     x1757            :in std_logic;
     x1758            :in std_logic;
     x1759            :in std_logic;
     x1760            :in std_logic;
     x1761            :in std_logic;
     x1762            :in std_logic;
     x1763            :in std_logic;
     x1764            :in std_logic;
     x1765            :in std_logic;
     x1766            :in std_logic;
     x1767            :in std_logic;
     x1768            :in std_logic;
     x1769            :in std_logic;
     x1770            :in std_logic;
     x1771            :in std_logic;
     x1772            :in std_logic;
     x1773            :in std_logic;
     x1774            :in std_logic;
     x1775            :in std_logic;
     x1776            :in std_logic;
     x1777            :in std_logic;
     x1778            :in std_logic;
     x1779            :in std_logic;
     x1780            :in std_logic;
     x1781            :in std_logic;
     x1782            :in std_logic;
     x1783            :in std_logic;
     x1784            :in std_logic;
     x1785            :in std_logic;
     x1786            :in std_logic;
     x1787            :in std_logic;
     x1788            :in std_logic;
     x1789            :in std_logic;
     x1790            :in std_logic;
     x1791            :in std_logic;
     x1792            :in std_logic;
     x1793            :in std_logic;
     x1794            :in std_logic;
     x1795            :in std_logic;
     x1796            :in std_logic;
     x1797            :in std_logic;
     x1798            :in std_logic;
     x1799            :in std_logic;
     x1800            :in std_logic;
     x1801            :in std_logic;
     x1802            :in std_logic;
     x1803            :in std_logic;
     x1804            :in std_logic;
     x1805            :in std_logic;
     x1806            :in std_logic;
     x1807            :in std_logic;
     x1808            :in std_logic;
     x1809            :in std_logic;
     x1810            :in std_logic;
     x1811            :in std_logic;
     x1812            :in std_logic;
     x1813            :in std_logic;
     x1814            :in std_logic;
     x1815            :in std_logic;
     x1816            :in std_logic;
     x1817            :in std_logic;
     x1818            :in std_logic;
     x1819            :in std_logic;
     x1820            :in std_logic;
     x1821            :in std_logic;
     x1822            :in std_logic;
     x1823            :in std_logic;
     x1824            :in std_logic;
     x1825            :in std_logic;
     x1826            :in std_logic;
     x1827            :in std_logic;
     x1828            :in std_logic;
     x1829            :in std_logic;
     x1830            :in std_logic;
     x1831            :in std_logic;
     x1832            :in std_logic;
     x1833            :in std_logic;
     x1834            :in std_logic;
     x1835            :in std_logic;
     x1836            :in std_logic;
     x1837            :in std_logic;
     x1838            :in std_logic;
     x1839            :in std_logic;
     x1840            :in std_logic;
     x1841            :in std_logic;
     x1842            :in std_logic;
     x1843            :in std_logic;
     x1844            :in std_logic;
     x1845            :in std_logic;
     x1846            :in std_logic;
     x1847            :in std_logic;
     x1848            :in std_logic;
     x1849            :in std_logic;
     x1850            :in std_logic;
     x1851            :in std_logic;
     x1852            :in std_logic;
     x1853            :in std_logic;
     x1854            :in std_logic;
     x1855            :in std_logic;
     x1856            :in std_logic;
     x1857            :in std_logic;
     x1858            :in std_logic;
     x1859            :in std_logic;
     x1860            :in std_logic;
     x1861            :in std_logic;
     x1862            :in std_logic;
     x1863            :in std_logic;
     x1864            :in std_logic;
     x1865            :in std_logic;
     x1866            :in std_logic;
     x1867            :in std_logic;
     x1868            :in std_logic;
     x1869            :in std_logic;
     x1870            :in std_logic;
     x1871            :in std_logic;
     x1872            :in std_logic;
     x1873            :in std_logic;
     x1874            :in std_logic;
     x1875            :in std_logic;
     x1876            :in std_logic;
     x1877            :in std_logic;
     x1878            :in std_logic;
     x1879            :in std_logic;
     x1880            :in std_logic;
     x1881            :in std_logic;
     x1882            :in std_logic;
     x1883            :in std_logic;
     x1884            :in std_logic;
     x1885            :in std_logic;
     x1886            :in std_logic;
     x1887            :in std_logic;
     x1888            :in std_logic;
     x1889            :in std_logic;
     x1890            :in std_logic;
     x1891            :in std_logic;
     x1892            :in std_logic;
     x1893            :in std_logic;
     x1894            :in std_logic;
     x1895            :in std_logic;
     x1896            :in std_logic;
     x1897            :in std_logic;
     x1898            :in std_logic;
     x1899            :in std_logic;
     x1900            :in std_logic;
     x1901            :in std_logic;
     x1902            :in std_logic;
     x1903            :in std_logic;
     x1904            :in std_logic;
     x1905            :in std_logic;
     x1906            :in std_logic;
     x1907            :in std_logic;
     x1908            :in std_logic;
     x1909            :in std_logic;
     x1910            :in std_logic;
     x1911            :in std_logic;
     x1912            :in std_logic;
     x1913            :in std_logic;
     x1914            :in std_logic;
     x1915            :in std_logic;
     x1916            :in std_logic;
     x1917            :in std_logic;
     x1918            :in std_logic;
     x1919            :in std_logic;
     x1920            :in std_logic;
     x1921            :in std_logic;
     x1922            :in std_logic;
     x1923            :in std_logic;
     x1924            :in std_logic;
     x1925            :in std_logic;
     x1926            :in std_logic;
     x1927            :in std_logic;
     x1928            :in std_logic;
     x1929            :in std_logic;
     x1930            :in std_logic;
     x1931            :in std_logic;
     x1932            :in std_logic;
     x1933            :in std_logic;
     x1934            :in std_logic;
     x1935            :in std_logic;
     x1936            :in std_logic;
     x1937            :in std_logic;
     x1938            :in std_logic;
     x1939            :in std_logic;
     x1940            :in std_logic;
     x1941            :in std_logic;
     x1942            :in std_logic;
     x1943            :in std_logic;
     x1944            :in std_logic;
     x1945            :in std_logic;
     x1946            :in std_logic;
     x1947            :in std_logic;
     x1948            :in std_logic;
     x1949            :in std_logic;
     x1950            :in std_logic;
     x1951            :in std_logic;
     x1952            :in std_logic;
     x1953            :in std_logic;
     x1954            :in std_logic;
     x1955            :in std_logic;
     x1956            :in std_logic;
     x1957            :in std_logic;
     x1958            :in std_logic;
     x1959            :in std_logic;
     x1960            :in std_logic;
     x1961            :in std_logic;
     x1962            :in std_logic;
     x1963            :in std_logic;
     x1964            :in std_logic;
     x1965            :in std_logic;
     x1966            :in std_logic;
     x1967            :in std_logic;
     x1968            :in std_logic;
     x1969            :in std_logic;
     x1970            :in std_logic;
     x1971            :in std_logic;
     x1972            :in std_logic;
     x1973            :in std_logic;
     x1974            :in std_logic;
     x1975            :in std_logic;
     x1976            :in std_logic;
     x1977            :in std_logic;
     x1978            :in std_logic;
     x1979            :in std_logic;
     x1980            :in std_logic;
     x1981            :in std_logic;
     x1982            :in std_logic;
     x1983            :in std_logic;
     x1984            :in std_logic;
     x1985            :in std_logic;
     x1986            :in std_logic;
     x1987            :in std_logic;
     x1988            :in std_logic;
     x1989            :in std_logic;
     x1990            :in std_logic;
     x1991            :in std_logic;
     x1992            :in std_logic;
     x1993            :in std_logic;
     x1994            :in std_logic;
     x1995            :in std_logic;
     x1996            :in std_logic;
     x1997            :in std_logic;
     x1998            :in std_logic;
     x1999            :in std_logic;
     x2000            :in std_logic;
     x2001            :in std_logic;
     x2002            :in std_logic;
     x2003            :in std_logic;
     x2004            :in std_logic;
     x2005            :in std_logic;
     x2006            :in std_logic;
     x2007            :in std_logic;
     x2008            :in std_logic;
     x2009            :in std_logic;
     x2010            :in std_logic;
     x2011            :in std_logic;
     x2012            :in std_logic;
     x2013            :in std_logic;
     x2014            :in std_logic;
     x2015            :in std_logic;
     x2016            :in std_logic;
     x2017            :in std_logic;
     x2018            :in std_logic;
     x2019            :in std_logic;
     x2020            :in std_logic;
     x2021            :in std_logic;
     x2022            :in std_logic;
     x2023            :in std_logic;
     x2024            :in std_logic;
     x2025            :in std_logic;
     x2026            :in std_logic;
     x2027            :in std_logic;
     x2028            :in std_logic;
     x2029            :in std_logic;
     x2030            :in std_logic;
     x2031            :in std_logic;
     x2032            :in std_logic;
     x2033            :in std_logic;
     x2034            :in std_logic;
     x2035            :in std_logic;
     x2036            :in std_logic;
     x2037            :in std_logic;
     x2038            :in std_logic;
     x2039            :in std_logic;
     x2040            :in std_logic;
     x2041            :in std_logic;
     x2042            :in std_logic;
     x2043            :in std_logic;
     x2044            :in std_logic;
     x2045            :in std_logic;
     x2046            :in std_logic;
     x2047            :in std_logic;
     x2048            :in std_logic;
     x2049            :in std_logic;
     x2050            :in std_logic;
     x2051            :in std_logic;
     x2052            :in std_logic;
     x2053            :in std_logic;
     x2054            :in std_logic;
     x2055            :in std_logic;
     x2056            :in std_logic;
     x2057            :in std_logic;
     x2058            :in std_logic;
     x2059            :in std_logic;
     x2060            :in std_logic;
     x2061            :in std_logic;
     x2062            :in std_logic;
     x2063            :in std_logic;
     x2064            :in std_logic;
     x2065            :in std_logic;
     x2066            :in std_logic;
     x2067            :in std_logic;
     x2068            :in std_logic;
     x2069            :in std_logic;
     x2070            :in std_logic;
     x2071            :in std_logic;
     x2072            :in std_logic;
     x2073            :in std_logic;
     x2074            :in std_logic;
     x2075            :in std_logic;
     x2076            :in std_logic;
     x2077            :in std_logic;
     x2078            :in std_logic;
     x2079            :in std_logic;
     x2080            :in std_logic;
     x2081            :in std_logic;
     x2082            :in std_logic;
     x2083            :in std_logic;
     x2084            :in std_logic;
     x2085            :in std_logic;
     x2086            :in std_logic;
     x2087            :in std_logic;
     x2088            :in std_logic;
     x2089            :in std_logic;
     x2090            :in std_logic;
     x2091            :in std_logic;
     x2092            :in std_logic;
     x2093            :in std_logic;
     x2094            :in std_logic;
     x2095            :in std_logic;
     x2096            :in std_logic;
     x2097            :in std_logic;
     x2098            :in std_logic;
     x2099            :in std_logic;
     x2100            :in std_logic;
     x2101            :in std_logic;
     x2102            :in std_logic;
     x2103            :in std_logic;
     x2104            :in std_logic;
     x2105            :in std_logic;
     x2106            :in std_logic;
     x2107            :in std_logic;
     x2108            :in std_logic;
     x2109            :in std_logic;
     x2110            :in std_logic;
     x2111            :in std_logic;
     x2112            :in std_logic;
     x2113            :in std_logic;
     x2114            :in std_logic;
     x2115            :in std_logic;
     x2116            :in std_logic;
     x2117            :in std_logic;
     x2118            :in std_logic;
     x2119            :in std_logic;
     x2120            :in std_logic;
     x2121            :in std_logic;
     x2122            :in std_logic;
     x2123            :in std_logic;
     x2124            :in std_logic;
     x2125            :in std_logic;
     x2126            :in std_logic;
     x2127            :in std_logic;
     x2128            :in std_logic;
     x2129            :in std_logic;
     x2130            :in std_logic;
     x2131            :in std_logic;
     x2132            :in std_logic;
     x2133            :in std_logic;
     x2134            :in std_logic;
     x2135            :in std_logic;
     x2136            :in std_logic;
     x2137            :in std_logic;
     x2138            :in std_logic;
     x2139            :in std_logic;
     x2140            :in std_logic;
     x2141            :in std_logic;
     x2142            :in std_logic;
     x2143            :in std_logic;
     x2144            :in std_logic;
     x2145            :in std_logic;
     x2146            :in std_logic;
     x2147            :in std_logic;
     x2148            :in std_logic;
     x2149            :in std_logic;
     x2150            :in std_logic;
     x2151            :in std_logic;
     x2152            :in std_logic;
     x2153            :in std_logic;
     x2154            :in std_logic;
     x2155            :in std_logic;
     x2156            :in std_logic;
     x2157            :in std_logic;
     x2158            :in std_logic;
     x2159            :in std_logic;
     x2160            :in std_logic;
     x2161            :in std_logic;
     x2162            :in std_logic;
     x2163            :in std_logic;
     x2164            :in std_logic;
     x2165            :in std_logic;
     x2166            :in std_logic;
     x2167            :in std_logic;
     x2168            :in std_logic;
     x2169            :in std_logic;
     x2170            :in std_logic;
     x2171            :in std_logic;
     x2172            :in std_logic;
     x2173            :in std_logic;
     x2174            :in std_logic;
     x2175            :in std_logic;
     x2176            :in std_logic;
     x2177            :in std_logic;
     x2178            :in std_logic;
     x2179            :in std_logic;
     x2180            :in std_logic;
     x2181            :in std_logic;
     x2182            :in std_logic;
     x2183            :in std_logic;
     x2184            :in std_logic;
     x2185            :in std_logic;
     x2186            :in std_logic;
     x2187            :in std_logic;
     x2188            :in std_logic;
     x2189            :in std_logic;
     x2190            :in std_logic;
     x2191            :in std_logic;
     x2192            :in std_logic;
     x2193            :in std_logic;
     x2194            :in std_logic;
     x2195            :in std_logic;
     x2196            :in std_logic;
     x2197            :in std_logic;
     x2198            :in std_logic;
     x2199            :in std_logic;
     x2200            :in std_logic;
     x2201            :in std_logic;
     x2202            :in std_logic;
     x2203            :in std_logic;
     x2204            :in std_logic;
     x2205            :in std_logic;
     x2206            :in std_logic;
     x2207            :in std_logic;
     x2208            :in std_logic;
     x2209            :in std_logic;
     x2210            :in std_logic;
     x2211            :in std_logic;
     x2212            :in std_logic;
     x2213            :in std_logic;
     x2214            :in std_logic;
     x2215            :in std_logic;
     x2216            :in std_logic;
     x2217            :in std_logic;
     x2218            :in std_logic;
     x2219            :in std_logic;
     x2220            :in std_logic;
     x2221            :in std_logic;
     x2222            :in std_logic;
     x2223            :in std_logic;
     x2224            :in std_logic;
     x2225            :in std_logic;
     x2226            :in std_logic;
     x2227            :in std_logic;
     x2228            :in std_logic;
     x2229            :in std_logic;
     x2230            :in std_logic;
     x2231            :in std_logic;
     x2232            :in std_logic;
     x2233            :in std_logic;
     x2234            :in std_logic;
     x2235            :in std_logic;
     x2236            :in std_logic;
     x2237            :in std_logic;
     x2238            :in std_logic;
     x2239            :in std_logic;
     x2240            :in std_logic;
     x2241            :in std_logic;
     x2242            :in std_logic;
     x2243            :in std_logic;
     x2244            :in std_logic;
     x2245            :in std_logic;
     x2246            :in std_logic;
     x2247            :in std_logic;
     x2248            :in std_logic;
     x2249            :in std_logic;
     x2250            :in std_logic;
     x2251            :in std_logic;
     x2252            :in std_logic;
     x2253            :in std_logic;
     x2254            :in std_logic;
     x2255            :in std_logic;
     x2256            :in std_logic;
     x2257            :in std_logic;
     x2258            :in std_logic;
     x2259            :in std_logic;
     x2260            :in std_logic;
     x2261            :in std_logic;
     x2262            :in std_logic;
     x2263            :in std_logic;
     x2264            :in std_logic;
     x2265            :in std_logic;
     x2266            :in std_logic;
     x2267            :in std_logic;
     x2268            :in std_logic;
     x2269            :in std_logic;
     x2270            :in std_logic;
     x2271            :in std_logic;
     x2272            :in std_logic;
     x2273            :in std_logic;
     x2274            :in std_logic;
     x2275            :in std_logic;
     x2276            :in std_logic;
     x2277            :in std_logic;
     x2278            :in std_logic;
     x2279            :in std_logic;
     x2280            :in std_logic;
     x2281            :in std_logic;
     x2282            :in std_logic;
     x2283            :in std_logic;
     x2284            :in std_logic;
     x2285            :in std_logic;
     x2286            :in std_logic;
     x2287            :in std_logic;
     x2288            :in std_logic;
     x2289            :in std_logic;
     x2290            :in std_logic;
     x2291            :in std_logic;
     x2292            :in std_logic;
     x2293            :in std_logic;
     x2294            :in std_logic;
     x2295            :in std_logic;
     x2296            :in std_logic;
     x2297            :in std_logic;
     x2298            :in std_logic;
     x2299            :in std_logic;
     x2300            :in std_logic;
     x2301            :in std_logic;
     x2302            :in std_logic;
     x2303            :in std_logic;
     x2304            :in std_logic;
     nbr_iter       : out std_logic_vector(4 downto 0);
     end_decision   :out std_logic
);
END component;

component FSM is
port ( clk, rst, start   : in std_logic;
stop_vnpu, stop_cnpu, stop_dec     : in std_logic;
start_vnpu, start_cnpu, start_decision : out std_logic;
end_decode         : out std_logic;
cpt_decision         : in std_logic_vector(2 downto 0));
end component;

FOR ALL : FSM
   USE ENTITY work.FSM(arch);
FOR ALL : decision
   USE ENTITY work.decision(arch_decision);
FOR ALL : ldpc
   USE ENTITY work.ldpc(ldpc_arch);

----------------------------- Declaration des Signaux -------------------
 signal s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,s958,s959,s960,s961,s962,s963,s964,s965,s966,s967,s968,s969,s970,s971,s972,s973,s974,s975,s976,s977,s978,s979,s980,s981,s982,s983,s984,s985,s986,s987,s988,s989,s990,s991,s992,s993,s994,s995,s996,s997,s998,s999,s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032,s1033,s1034,s1035,s1036,s1037,s1038,s1039,s1040,s1041,s1042,s1043,s1044,s1045,s1046,s1047,s1048,s1049,s1050,s1051,s1052,s1053,s1054,s1055,s1056,s1057,s1058,s1059,s1060,s1061,s1062,s1063,s1064,s1065,s1066,s1067,s1068,s1069,s1070,s1071,s1072,s1073,s1074,s1075,s1076,s1077,s1078,s1079,s1080,s1081,s1082,s1083,s1084,s1085,s1086,s1087,s1088,s1089,s1090,s1091,s1092,s1093,s1094,s1095,s1096,s1097,s1098,s1099,s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124,s1125,s1126,s1127,s1128,s1129,s1130,s1131,s1132,s1133,s1134,s1135,s1136,s1137,s1138,s1139,s1140,s1141,s1142,s1143,s1144,s1145,s1146,s1147,s1148,s1149,s1150,s1151,s1152,s1153,s1154,s1155,s1156,s1157,s1158,s1159,s1160,s1161,s1162,s1163,s1164,s1165,s1166,s1167,s1168,s1169,s1170,s1171,s1172,s1173,s1174,s1175,s1176,s1177,s1178,s1179,s1180,s1181,s1182,s1183,s1184,s1185,s1186,s1187,s1188,s1189,s1190,s1191,s1192,s1193,s1194,s1195,s1196,s1197,s1198,s1199,s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,s1231,s1232,s1233,s1234,s1235,s1236,s1237,s1238,s1239,s1240,s1241,s1242,s1243,s1244,s1245,s1246,s1247,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255,s1256,s1257,s1258,s1259,s1260,s1261,s1262,s1263,s1264,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272,s1273,s1274,s1275,s1276,s1277,s1278,s1279,s1280,s1281,s1282,s1283,s1284,s1285,s1286,s1287,s1288,s1289,s1290,s1291,s1292,s1293,s1294,s1295,s1296,s1297,s1298,s1299,s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324,s1325,s1326,s1327,s1328,s1329,s1330,s1331,s1332,s1333,s1334,s1335,s1336,s1337,s1338,s1339,s1340,s1341,s1342,s1343,s1344,s1345,s1346,s1347,s1348,s1349,s1350,s1351,s1352,s1353,s1354,s1355,s1356,s1357,s1358,s1359,s1360,s1361,s1362,s1363,s1364,s1365,s1366,s1367,s1368,s1369,s1370,s1371,s1372,s1373,s1374,s1375,s1376,s1377,s1378,s1379,s1380,s1381,s1382,s1383,s1384,s1385,s1386,s1387,s1388,s1389,s1390,s1391,s1392,s1393,s1394,s1395,s1396,s1397,s1398,s1399,s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425,s1426,s1427,s1428,s1429,s1430,s1431,s1432,s1433,s1434,s1435,s1436,s1437,s1438,s1439,s1440,s1441,s1442,s1443,s1444,s1445,s1446,s1447,s1448,s1449,s1450,s1451,s1452,s1453,s1454,s1455,s1456,s1457,s1458,s1459,s1460,s1461,s1462,s1463,s1464,s1465,s1466,s1467,s1468,s1469,s1470,s1471,s1472,s1473,s1474,s1475,s1476,s1477,s1478,s1479,s1480,s1481,s1482,s1483,s1484,s1485,s1486,s1487,s1488,s1489,s1490,s1491,s1492,s1493,s1494,s1495,s1496,s1497,s1498,s1499,s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,s1520,s1521,s1522,s1523,s1524,s1525,s1526,s1527,s1528,s1529,s1530,s1531,s1532,s1533,s1534,s1535,s1536,s1537,s1538,s1539,s1540,s1541,s1542,s1543,s1544,s1545,s1546,s1547,s1548,s1549,s1550,s1551,s1552,s1553,s1554,s1555,s1556,s1557,s1558,s1559,s1560,s1561,s1562,s1563,s1564,s1565,s1566,s1567,s1568,s1569,s1570,s1571,s1572,s1573,s1574,s1575,s1576,s1577,s1578,s1579,s1580,s1581,s1582,s1583,s1584,s1585,s1586,s1587,s1588,s1589,s1590,s1591,s1592,s1593,s1594,s1595,s1596,s1597,s1598,s1599,s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624,s1625,s1626,s1627,s1628,s1629,s1630,s1631,s1632,s1633,s1634,s1635,s1636,s1637,s1638,s1639,s1640,s1641,s1642,s1643,s1644,s1645,s1646,s1647,s1648,s1649,s1650,s1651,s1652,s1653,s1654,s1655,s1656,s1657,s1658,s1659,s1660,s1661,s1662,s1663,s1664,s1665,s1666,s1667,s1668,s1669,s1670,s1671,s1672,s1673,s1674,s1675,s1676,s1677,s1678,s1679,s1680,s1681,s1682,s1683,s1684,s1685,s1686,s1687,s1688,s1689,s1690,s1691,s1692,s1693,s1694,s1695,s1696,s1697,s1698,s1699,s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724,s1725,s1726,s1727,s1728,s1729,s1730,s1731,s1732,s1733,s1734,s1735,s1736,s1737,s1738,s1739,s1740,s1741,s1742,s1743,s1744,s1745,s1746,s1747,s1748,s1749,s1750,s1751,s1752,s1753,s1754,s1755,s1756,s1757,s1758,s1759,s1760,s1761,s1762,s1763,s1764,s1765,s1766,s1767,s1768,s1769,s1770,s1771,s1772,s1773,s1774,s1775,s1776,s1777,s1778,s1779,s1780,s1781,s1782,s1783,s1784,s1785,s1786,s1787,s1788,s1789,s1790,s1791,s1792,s1793,s1794,s1795,s1796,s1797,s1798,s1799,s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824,s1825,s1826,s1827,s1828,s1829,s1830,s1831,s1832,s1833,s1834,s1835,s1836,s1837,s1838,s1839,s1840,s1841,s1842,s1843,s1844,s1845,s1846,s1847,s1848,s1849,s1850,s1851,s1852,s1853,s1854,s1855,s1856,s1857,s1858,s1859,s1860,s1861,s1862,s1863,s1864,s1865,s1866,s1867,s1868,s1869,s1870,s1871,s1872,s1873,s1874,s1875,s1876,s1877,s1878,s1879,s1880,s1881,s1882,s1883,s1884,s1885,s1886,s1887,s1888,s1889,s1890,s1891,s1892,s1893,s1894,s1895,s1896,s1897,s1898,s1899,s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,s1920,s1921,s1922,s1923,s1924,s1925,s1926,s1927,s1928,s1929,s1930,s1931,s1932,s1933,s1934,s1935,s1936,s1937,s1938,s1939,s1940,s1941,s1942,s1943,s1944,s1945,s1946,s1947,s1948,s1949,s1950,s1951,s1952,s1953,s1954,s1955,s1956,s1957,s1958,s1959,s1960,s1961,s1962,s1963,s1964,s1965,s1966,s1967,s1968,s1969,s1970,s1971,s1972,s1973,s1974,s1975,s1976,s1977,s1978,s1979,s1980,s1981,s1982,s1983,s1984,s1985,s1986,s1987,s1988,s1989,s1990,s1991,s1992,s1993,s1994,s1995,s1996,s1997,s1998,s1999,s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024,s2025,s2026,s2027,s2028,s2029,s2030,s2031,s2032,s2033,s2034,s2035,s2036,s2037,s2038,s2039,s2040,s2041,s2042,s2043,s2044,s2045,s2046,s2047,s2048,s2049,s2050,s2051,s2052,s2053,s2054,s2055,s2056,s2057,s2058,s2059,s2060,s2061,s2062,s2063,s2064,s2065,s2066,s2067,s2068,s2069,s2070,s2071,s2072,s2073,s2074,s2075,s2076,s2077,s2078,s2079,s2080,s2081,s2082,s2083,s2084,s2085,s2086,s2087,s2088,s2089,s2090,s2091,s2092,s2093,s2094,s2095,s2096,s2097,s2098,s2099,s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124,s2125,s2126,s2127,s2128,s2129,s2130,s2131,s2132,s2133,s2134,s2135,s2136,s2137,s2138,s2139,s2140,s2141,s2142,s2143,s2144,s2145,s2146,s2147,s2148,s2149,s2150,s2151,s2152,s2153,s2154,s2155,s2156,s2157,s2158,s2159,s2160,s2161,s2162,s2163,s2164,s2165,s2166,s2167,s2168,s2169,s2170,s2171,s2172,s2173,s2174,s2175,s2176,s2177,s2178,s2179,s2180,s2181,s2182,s2183,s2184,s2185,s2186,s2187,s2188,s2189,s2190,s2191,s2192,s2193,s2194,s2195,s2196,s2197,s2198,s2199,s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224,s2225,s2226,s2227,s2228,s2229,s2230,s2231,s2232,s2233,s2234,s2235,s2236,s2237,s2238,s2239,s2240,s2241,s2242,s2243,s2244,s2245,s2246,s2247,s2248,s2249,s2250,s2251,s2252,s2253,s2254,s2255,s2256,s2257,s2258,s2259,s2260,s2261,s2262,s2263,s2264,s2265,s2266,s2267,s2268,s2269,s2270,s2271,s2272,s2273,s2274,s2275,s2276,s2277,s2278,s2279,s2280,s2281,s2282,s2283,s2284,s2285,s2286,s2287,s2288,s2289,s2290,s2291,s2292,s2293,s2294,s2295,s2296,s2297,s2298,s2299,s2300,s2301,s2302,s2303,s2304:std_logic;
SIGNAL x_x,y_y,startcn,startvn           :std_logic;
SIGNAL str_parity,stop_de                 : std_logic;
signal ctc                                : std_logic_vector(2 downto 0):="111";

begin
----------------------------- maping les components -------------------
 FSM1:FSM
port map (
     clk=>clock,
	  rst=>reset,
	  start=>start_decoder,
	  stop_cnpu=> x_x,
	  stop_vnpu=> y_y,
	  stop_dec=>stop_de,
	  start_cnpu=>startcn,
	  start_vnpu=>startvn,
	  start_decision=>str_parity,
	  end_decode=>end_decoder,
   	  cpt_decision=>ctc
       );

decision1:decision port map(clock,reset,str_parity,iter_Mx,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,s958,s959,s960,s961,s962,s963,s964,s965,s966,s967,s968,s969,s970,s971,s972,s973,s974,s975,s976,s977,s978,s979,s980,s981,s982,s983,s984,s985,s986,s987,s988,s989,s990,s991,s992,s993,s994,s995,s996,s997,s998,s999,s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032,s1033,s1034,s1035,s1036,s1037,s1038,s1039,s1040,s1041,s1042,s1043,s1044,s1045,s1046,s1047,s1048,s1049,s1050,s1051,s1052,s1053,s1054,s1055,s1056,s1057,s1058,s1059,s1060,s1061,s1062,s1063,s1064,s1065,s1066,s1067,s1068,s1069,s1070,s1071,s1072,s1073,s1074,s1075,s1076,s1077,s1078,s1079,s1080,s1081,s1082,s1083,s1084,s1085,s1086,s1087,s1088,s1089,s1090,s1091,s1092,s1093,s1094,s1095,s1096,s1097,s1098,s1099,s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124,s1125,s1126,s1127,s1128,s1129,s1130,s1131,s1132,s1133,s1134,s1135,s1136,s1137,s1138,s1139,s1140,s1141,s1142,s1143,s1144,s1145,s1146,s1147,s1148,s1149,s1150,s1151,s1152,s1153,s1154,s1155,s1156,s1157,s1158,s1159,s1160,s1161,s1162,s1163,s1164,s1165,s1166,s1167,s1168,s1169,s1170,s1171,s1172,s1173,s1174,s1175,s1176,s1177,s1178,s1179,s1180,s1181,s1182,s1183,s1184,s1185,s1186,s1187,s1188,s1189,s1190,s1191,s1192,s1193,s1194,s1195,s1196,s1197,s1198,s1199,s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,s1231,s1232,s1233,s1234,s1235,s1236,s1237,s1238,s1239,s1240,s1241,s1242,s1243,s1244,s1245,s1246,s1247,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255,s1256,s1257,s1258,s1259,s1260,s1261,s1262,s1263,s1264,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272,s1273,s1274,s1275,s1276,s1277,s1278,s1279,s1280,s1281,s1282,s1283,s1284,s1285,s1286,s1287,s1288,s1289,s1290,s1291,s1292,s1293,s1294,s1295,s1296,s1297,s1298,s1299,s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324,s1325,s1326,s1327,s1328,s1329,s1330,s1331,s1332,s1333,s1334,s1335,s1336,s1337,s1338,s1339,s1340,s1341,s1342,s1343,s1344,s1345,s1346,s1347,s1348,s1349,s1350,s1351,s1352,s1353,s1354,s1355,s1356,s1357,s1358,s1359,s1360,s1361,s1362,s1363,s1364,s1365,s1366,s1367,s1368,s1369,s1370,s1371,s1372,s1373,s1374,s1375,s1376,s1377,s1378,s1379,s1380,s1381,s1382,s1383,s1384,s1385,s1386,s1387,s1388,s1389,s1390,s1391,s1392,s1393,s1394,s1395,s1396,s1397,s1398,s1399,s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425,s1426,s1427,s1428,s1429,s1430,s1431,s1432,s1433,s1434,s1435,s1436,s1437,s1438,s1439,s1440,s1441,s1442,s1443,s1444,s1445,s1446,s1447,s1448,s1449,s1450,s1451,s1452,s1453,s1454,s1455,s1456,s1457,s1458,s1459,s1460,s1461,s1462,s1463,s1464,s1465,s1466,s1467,s1468,s1469,s1470,s1471,s1472,s1473,s1474,s1475,s1476,s1477,s1478,s1479,s1480,s1481,s1482,s1483,s1484,s1485,s1486,s1487,s1488,s1489,s1490,s1491,s1492,s1493,s1494,s1495,s1496,s1497,s1498,s1499,s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,s1520,s1521,s1522,s1523,s1524,s1525,s1526,s1527,s1528,s1529,s1530,s1531,s1532,s1533,s1534,s1535,s1536,s1537,s1538,s1539,s1540,s1541,s1542,s1543,s1544,s1545,s1546,s1547,s1548,s1549,s1550,s1551,s1552,s1553,s1554,s1555,s1556,s1557,s1558,s1559,s1560,s1561,s1562,s1563,s1564,s1565,s1566,s1567,s1568,s1569,s1570,s1571,s1572,s1573,s1574,s1575,s1576,s1577,s1578,s1579,s1580,s1581,s1582,s1583,s1584,s1585,s1586,s1587,s1588,s1589,s1590,s1591,s1592,s1593,s1594,s1595,s1596,s1597,s1598,s1599,s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624,s1625,s1626,s1627,s1628,s1629,s1630,s1631,s1632,s1633,s1634,s1635,s1636,s1637,s1638,s1639,s1640,s1641,s1642,s1643,s1644,s1645,s1646,s1647,s1648,s1649,s1650,s1651,s1652,s1653,s1654,s1655,s1656,s1657,s1658,s1659,s1660,s1661,s1662,s1663,s1664,s1665,s1666,s1667,s1668,s1669,s1670,s1671,s1672,s1673,s1674,s1675,s1676,s1677,s1678,s1679,s1680,s1681,s1682,s1683,s1684,s1685,s1686,s1687,s1688,s1689,s1690,s1691,s1692,s1693,s1694,s1695,s1696,s1697,s1698,s1699,s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724,s1725,s1726,s1727,s1728,s1729,s1730,s1731,s1732,s1733,s1734,s1735,s1736,s1737,s1738,s1739,s1740,s1741,s1742,s1743,s1744,s1745,s1746,s1747,s1748,s1749,s1750,s1751,s1752,s1753,s1754,s1755,s1756,s1757,s1758,s1759,s1760,s1761,s1762,s1763,s1764,s1765,s1766,s1767,s1768,s1769,s1770,s1771,s1772,s1773,s1774,s1775,s1776,s1777,s1778,s1779,s1780,s1781,s1782,s1783,s1784,s1785,s1786,s1787,s1788,s1789,s1790,s1791,s1792,s1793,s1794,s1795,s1796,s1797,s1798,s1799,s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824,s1825,s1826,s1827,s1828,s1829,s1830,s1831,s1832,s1833,s1834,s1835,s1836,s1837,s1838,s1839,s1840,s1841,s1842,s1843,s1844,s1845,s1846,s1847,s1848,s1849,s1850,s1851,s1852,s1853,s1854,s1855,s1856,s1857,s1858,s1859,s1860,s1861,s1862,s1863,s1864,s1865,s1866,s1867,s1868,s1869,s1870,s1871,s1872,s1873,s1874,s1875,s1876,s1877,s1878,s1879,s1880,s1881,s1882,s1883,s1884,s1885,s1886,s1887,s1888,s1889,s1890,s1891,s1892,s1893,s1894,s1895,s1896,s1897,s1898,s1899,s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,s1920,s1921,s1922,s1923,s1924,s1925,s1926,s1927,s1928,s1929,s1930,s1931,s1932,s1933,s1934,s1935,s1936,s1937,s1938,s1939,s1940,s1941,s1942,s1943,s1944,s1945,s1946,s1947,s1948,s1949,s1950,s1951,s1952,s1953,s1954,s1955,s1956,s1957,s1958,s1959,s1960,s1961,s1962,s1963,s1964,s1965,s1966,s1967,s1968,s1969,s1970,s1971,s1972,s1973,s1974,s1975,s1976,s1977,s1978,s1979,s1980,s1981,s1982,s1983,s1984,s1985,s1986,s1987,s1988,s1989,s1990,s1991,s1992,s1993,s1994,s1995,s1996,s1997,s1998,s1999,s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024,s2025,s2026,s2027,s2028,s2029,s2030,s2031,s2032,s2033,s2034,s2035,s2036,s2037,s2038,s2039,s2040,s2041,s2042,s2043,s2044,s2045,s2046,s2047,s2048,s2049,s2050,s2051,s2052,s2053,s2054,s2055,s2056,s2057,s2058,s2059,s2060,s2061,s2062,s2063,s2064,s2065,s2066,s2067,s2068,s2069,s2070,s2071,s2072,s2073,s2074,s2075,s2076,s2077,s2078,s2079,s2080,s2081,s2082,s2083,s2084,s2085,s2086,s2087,s2088,s2089,s2090,s2091,s2092,s2093,s2094,s2095,s2096,s2097,s2098,s2099,s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124,s2125,s2126,s2127,s2128,s2129,s2130,s2131,s2132,s2133,s2134,s2135,s2136,s2137,s2138,s2139,s2140,s2141,s2142,s2143,s2144,s2145,s2146,s2147,s2148,s2149,s2150,s2151,s2152,s2153,s2154,s2155,s2156,s2157,s2158,s2159,s2160,s2161,s2162,s2163,s2164,s2165,s2166,s2167,s2168,s2169,s2170,s2171,s2172,s2173,s2174,s2175,s2176,s2177,s2178,s2179,s2180,s2181,s2182,s2183,s2184,s2185,s2186,s2187,s2188,s2189,s2190,s2191,s2192,s2193,s2194,s2195,s2196,s2197,s2198,s2199,s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224,s2225,s2226,s2227,s2228,s2229,s2230,s2231,s2232,s2233,s2234,s2235,s2236,s2237,s2238,s2239,s2240,s2241,s2242,s2243,s2244,s2245,s2246,s2247,s2248,s2249,s2250,s2251,s2252,s2253,s2254,s2255,s2256,s2257,s2258,s2259,s2260,s2261,s2262,s2263,s2264,s2265,s2266,s2267,s2268,s2269,s2270,s2271,s2272,s2273,s2274,s2275,s2276,s2277,s2278,s2279,s2280,s2281,s2282,s2283,s2284,s2285,s2286,s2287,s2288,s2289,s2290,s2291,s2292,s2293,s2294,s2295,s2296,s2297,s2298,s2299,s2300,s2301,s2302,s2303,s2304,num_iter,stop_de);

ldpc1:ldpc port map(clock,reset,startvn,startcn,L1,L2,L3,L4,L5,L6,L7,L8,L9,L10,L11,L12,L13,L14,L15,L16,L17,L18,L19,L20,L21,L22,L23,L24,L25,L26,L27,L28,L29,L30,L31,L32,L33,L34,L35,L36,L37,L38,L39,L40,L41,L42,L43,L44,L45,L46,L47,L48,L49,L50,L51,L52,L53,L54,L55,L56,L57,L58,L59,L60,L61,L62,L63,L64,L65,L66,L67,L68,L69,L70,L71,L72,L73,L74,L75,L76,L77,L78,L79,L80,L81,L82,L83,L84,L85,L86,L87,L88,L89,L90,L91,L92,L93,L94,L95,L96,L97,L98,L99,L100,L101,L102,L103,L104,L105,L106,L107,L108,L109,L110,L111,L112,L113,L114,L115,L116,L117,L118,L119,L120,L121,L122,L123,L124,L125,L126,L127,L128,L129,L130,L131,L132,L133,L134,L135,L136,L137,L138,L139,L140,L141,L142,L143,L144,L145,L146,L147,L148,L149,L150,L151,L152,L153,L154,L155,L156,L157,L158,L159,L160,L161,L162,L163,L164,L165,L166,L167,L168,L169,L170,L171,L172,L173,L174,L175,L176,L177,L178,L179,L180,L181,L182,L183,L184,L185,L186,L187,L188,L189,L190,L191,L192,L193,L194,L195,L196,L197,L198,L199,L200,L201,L202,L203,L204,L205,L206,L207,L208,L209,L210,L211,L212,L213,L214,L215,L216,L217,L218,L219,L220,L221,L222,L223,L224,L225,L226,L227,L228,L229,L230,L231,L232,L233,L234,L235,L236,L237,L238,L239,L240,L241,L242,L243,L244,L245,L246,L247,L248,L249,L250,L251,L252,L253,L254,L255,L256,L257,L258,L259,L260,L261,L262,L263,L264,L265,L266,L267,L268,L269,L270,L271,L272,L273,L274,L275,L276,L277,L278,L279,L280,L281,L282,L283,L284,L285,L286,L287,L288,L289,L290,L291,L292,L293,L294,L295,L296,L297,L298,L299,L300,L301,L302,L303,L304,L305,L306,L307,L308,L309,L310,L311,L312,L313,L314,L315,L316,L317,L318,L319,L320,L321,L322,L323,L324,L325,L326,L327,L328,L329,L330,L331,L332,L333,L334,L335,L336,L337,L338,L339,L340,L341,L342,L343,L344,L345,L346,L347,L348,L349,L350,L351,L352,L353,L354,L355,L356,L357,L358,L359,L360,L361,L362,L363,L364,L365,L366,L367,L368,L369,L370,L371,L372,L373,L374,L375,L376,L377,L378,L379,L380,L381,L382,L383,L384,L385,L386,L387,L388,L389,L390,L391,L392,L393,L394,L395,L396,L397,L398,L399,L400,L401,L402,L403,L404,L405,L406,L407,L408,L409,L410,L411,L412,L413,L414,L415,L416,L417,L418,L419,L420,L421,L422,L423,L424,L425,L426,L427,L428,L429,L430,L431,L432,L433,L434,L435,L436,L437,L438,L439,L440,L441,L442,L443,L444,L445,L446,L447,L448,L449,L450,L451,L452,L453,L454,L455,L456,L457,L458,L459,L460,L461,L462,L463,L464,L465,L466,L467,L468,L469,L470,L471,L472,L473,L474,L475,L476,L477,L478,L479,L480,L481,L482,L483,L484,L485,L486,L487,L488,L489,L490,L491,L492,L493,L494,L495,L496,L497,L498,L499,L500,L501,L502,L503,L504,L505,L506,L507,L508,L509,L510,L511,L512,L513,L514,L515,L516,L517,L518,L519,L520,L521,L522,L523,L524,L525,L526,L527,L528,L529,L530,L531,L532,L533,L534,L535,L536,L537,L538,L539,L540,L541,L542,L543,L544,L545,L546,L547,L548,L549,L550,L551,L552,L553,L554,L555,L556,L557,L558,L559,L560,L561,L562,L563,L564,L565,L566,L567,L568,L569,L570,L571,L572,L573,L574,L575,L576,L577,L578,L579,L580,L581,L582,L583,L584,L585,L586,L587,L588,L589,L590,L591,L592,L593,L594,L595,L596,L597,L598,L599,L600,L601,L602,L603,L604,L605,L606,L607,L608,L609,L610,L611,L612,L613,L614,L615,L616,L617,L618,L619,L620,L621,L622,L623,L624,L625,L626,L627,L628,L629,L630,L631,L632,L633,L634,L635,L636,L637,L638,L639,L640,L641,L642,L643,L644,L645,L646,L647,L648,L649,L650,L651,L652,L653,L654,L655,L656,L657,L658,L659,L660,L661,L662,L663,L664,L665,L666,L667,L668,L669,L670,L671,L672,L673,L674,L675,L676,L677,L678,L679,L680,L681,L682,L683,L684,L685,L686,L687,L688,L689,L690,L691,L692,L693,L694,L695,L696,L697,L698,L699,L700,L701,L702,L703,L704,L705,L706,L707,L708,L709,L710,L711,L712,L713,L714,L715,L716,L717,L718,L719,L720,L721,L722,L723,L724,L725,L726,L727,L728,L729,L730,L731,L732,L733,L734,L735,L736,L737,L738,L739,L740,L741,L742,L743,L744,L745,L746,L747,L748,L749,L750,L751,L752,L753,L754,L755,L756,L757,L758,L759,L760,L761,L762,L763,L764,L765,L766,L767,L768,L769,L770,L771,L772,L773,L774,L775,L776,L777,L778,L779,L780,L781,L782,L783,L784,L785,L786,L787,L788,L789,L790,L791,L792,L793,L794,L795,L796,L797,L798,L799,L800,L801,L802,L803,L804,L805,L806,L807,L808,L809,L810,L811,L812,L813,L814,L815,L816,L817,L818,L819,L820,L821,L822,L823,L824,L825,L826,L827,L828,L829,L830,L831,L832,L833,L834,L835,L836,L837,L838,L839,L840,L841,L842,L843,L844,L845,L846,L847,L848,L849,L850,L851,L852,L853,L854,L855,L856,L857,L858,L859,L860,L861,L862,L863,L864,L865,L866,L867,L868,L869,L870,L871,L872,L873,L874,L875,L876,L877,L878,L879,L880,L881,L882,L883,L884,L885,L886,L887,L888,L889,L890,L891,L892,L893,L894,L895,L896,L897,L898,L899,L900,L901,L902,L903,L904,L905,L906,L907,L908,L909,L910,L911,L912,L913,L914,L915,L916,L917,L918,L919,L920,L921,L922,L923,L924,L925,L926,L927,L928,L929,L930,L931,L932,L933,L934,L935,L936,L937,L938,L939,L940,L941,L942,L943,L944,L945,L946,L947,L948,L949,L950,L951,L952,L953,L954,L955,L956,L957,L958,L959,L960,L961,L962,L963,L964,L965,L966,L967,L968,L969,L970,L971,L972,L973,L974,L975,L976,L977,L978,L979,L980,L981,L982,L983,L984,L985,L986,L987,L988,L989,L990,L991,L992,L993,L994,L995,L996,L997,L998,L999,L1000,L1001,L1002,L1003,L1004,L1005,L1006,L1007,L1008,L1009,L1010,L1011,L1012,L1013,L1014,L1015,L1016,L1017,L1018,L1019,L1020,L1021,L1022,L1023,L1024,L1025,L1026,L1027,L1028,L1029,L1030,L1031,L1032,L1033,L1034,L1035,L1036,L1037,L1038,L1039,L1040,L1041,L1042,L1043,L1044,L1045,L1046,L1047,L1048,L1049,L1050,L1051,L1052,L1053,L1054,L1055,L1056,L1057,L1058,L1059,L1060,L1061,L1062,L1063,L1064,L1065,L1066,L1067,L1068,L1069,L1070,L1071,L1072,L1073,L1074,L1075,L1076,L1077,L1078,L1079,L1080,L1081,L1082,L1083,L1084,L1085,L1086,L1087,L1088,L1089,L1090,L1091,L1092,L1093,L1094,L1095,L1096,L1097,L1098,L1099,L1100,L1101,L1102,L1103,L1104,L1105,L1106,L1107,L1108,L1109,L1110,L1111,L1112,L1113,L1114,L1115,L1116,L1117,L1118,L1119,L1120,L1121,L1122,L1123,L1124,L1125,L1126,L1127,L1128,L1129,L1130,L1131,L1132,L1133,L1134,L1135,L1136,L1137,L1138,L1139,L1140,L1141,L1142,L1143,L1144,L1145,L1146,L1147,L1148,L1149,L1150,L1151,L1152,L1153,L1154,L1155,L1156,L1157,L1158,L1159,L1160,L1161,L1162,L1163,L1164,L1165,L1166,L1167,L1168,L1169,L1170,L1171,L1172,L1173,L1174,L1175,L1176,L1177,L1178,L1179,L1180,L1181,L1182,L1183,L1184,L1185,L1186,L1187,L1188,L1189,L1190,L1191,L1192,L1193,L1194,L1195,L1196,L1197,L1198,L1199,L1200,L1201,L1202,L1203,L1204,L1205,L1206,L1207,L1208,L1209,L1210,L1211,L1212,L1213,L1214,L1215,L1216,L1217,L1218,L1219,L1220,L1221,L1222,L1223,L1224,L1225,L1226,L1227,L1228,L1229,L1230,L1231,L1232,L1233,L1234,L1235,L1236,L1237,L1238,L1239,L1240,L1241,L1242,L1243,L1244,L1245,L1246,L1247,L1248,L1249,L1250,L1251,L1252,L1253,L1254,L1255,L1256,L1257,L1258,L1259,L1260,L1261,L1262,L1263,L1264,L1265,L1266,L1267,L1268,L1269,L1270,L1271,L1272,L1273,L1274,L1275,L1276,L1277,L1278,L1279,L1280,L1281,L1282,L1283,L1284,L1285,L1286,L1287,L1288,L1289,L1290,L1291,L1292,L1293,L1294,L1295,L1296,L1297,L1298,L1299,L1300,L1301,L1302,L1303,L1304,L1305,L1306,L1307,L1308,L1309,L1310,L1311,L1312,L1313,L1314,L1315,L1316,L1317,L1318,L1319,L1320,L1321,L1322,L1323,L1324,L1325,L1326,L1327,L1328,L1329,L1330,L1331,L1332,L1333,L1334,L1335,L1336,L1337,L1338,L1339,L1340,L1341,L1342,L1343,L1344,L1345,L1346,L1347,L1348,L1349,L1350,L1351,L1352,L1353,L1354,L1355,L1356,L1357,L1358,L1359,L1360,L1361,L1362,L1363,L1364,L1365,L1366,L1367,L1368,L1369,L1370,L1371,L1372,L1373,L1374,L1375,L1376,L1377,L1378,L1379,L1380,L1381,L1382,L1383,L1384,L1385,L1386,L1387,L1388,L1389,L1390,L1391,L1392,L1393,L1394,L1395,L1396,L1397,L1398,L1399,L1400,L1401,L1402,L1403,L1404,L1405,L1406,L1407,L1408,L1409,L1410,L1411,L1412,L1413,L1414,L1415,L1416,L1417,L1418,L1419,L1420,L1421,L1422,L1423,L1424,L1425,L1426,L1427,L1428,L1429,L1430,L1431,L1432,L1433,L1434,L1435,L1436,L1437,L1438,L1439,L1440,L1441,L1442,L1443,L1444,L1445,L1446,L1447,L1448,L1449,L1450,L1451,L1452,L1453,L1454,L1455,L1456,L1457,L1458,L1459,L1460,L1461,L1462,L1463,L1464,L1465,L1466,L1467,L1468,L1469,L1470,L1471,L1472,L1473,L1474,L1475,L1476,L1477,L1478,L1479,L1480,L1481,L1482,L1483,L1484,L1485,L1486,L1487,L1488,L1489,L1490,L1491,L1492,L1493,L1494,L1495,L1496,L1497,L1498,L1499,L1500,L1501,L1502,L1503,L1504,L1505,L1506,L1507,L1508,L1509,L1510,L1511,L1512,L1513,L1514,L1515,L1516,L1517,L1518,L1519,L1520,L1521,L1522,L1523,L1524,L1525,L1526,L1527,L1528,L1529,L1530,L1531,L1532,L1533,L1534,L1535,L1536,L1537,L1538,L1539,L1540,L1541,L1542,L1543,L1544,L1545,L1546,L1547,L1548,L1549,L1550,L1551,L1552,L1553,L1554,L1555,L1556,L1557,L1558,L1559,L1560,L1561,L1562,L1563,L1564,L1565,L1566,L1567,L1568,L1569,L1570,L1571,L1572,L1573,L1574,L1575,L1576,L1577,L1578,L1579,L1580,L1581,L1582,L1583,L1584,L1585,L1586,L1587,L1588,L1589,L1590,L1591,L1592,L1593,L1594,L1595,L1596,L1597,L1598,L1599,L1600,L1601,L1602,L1603,L1604,L1605,L1606,L1607,L1608,L1609,L1610,L1611,L1612,L1613,L1614,L1615,L1616,L1617,L1618,L1619,L1620,L1621,L1622,L1623,L1624,L1625,L1626,L1627,L1628,L1629,L1630,L1631,L1632,L1633,L1634,L1635,L1636,L1637,L1638,L1639,L1640,L1641,L1642,L1643,L1644,L1645,L1646,L1647,L1648,L1649,L1650,L1651,L1652,L1653,L1654,L1655,L1656,L1657,L1658,L1659,L1660,L1661,L1662,L1663,L1664,L1665,L1666,L1667,L1668,L1669,L1670,L1671,L1672,L1673,L1674,L1675,L1676,L1677,L1678,L1679,L1680,L1681,L1682,L1683,L1684,L1685,L1686,L1687,L1688,L1689,L1690,L1691,L1692,L1693,L1694,L1695,L1696,L1697,L1698,L1699,L1700,L1701,L1702,L1703,L1704,L1705,L1706,L1707,L1708,L1709,L1710,L1711,L1712,L1713,L1714,L1715,L1716,L1717,L1718,L1719,L1720,L1721,L1722,L1723,L1724,L1725,L1726,L1727,L1728,L1729,L1730,L1731,L1732,L1733,L1734,L1735,L1736,L1737,L1738,L1739,L1740,L1741,L1742,L1743,L1744,L1745,L1746,L1747,L1748,L1749,L1750,L1751,L1752,L1753,L1754,L1755,L1756,L1757,L1758,L1759,L1760,L1761,L1762,L1763,L1764,L1765,L1766,L1767,L1768,L1769,L1770,L1771,L1772,L1773,L1774,L1775,L1776,L1777,L1778,L1779,L1780,L1781,L1782,L1783,L1784,L1785,L1786,L1787,L1788,L1789,L1790,L1791,L1792,L1793,L1794,L1795,L1796,L1797,L1798,L1799,L1800,L1801,L1802,L1803,L1804,L1805,L1806,L1807,L1808,L1809,L1810,L1811,L1812,L1813,L1814,L1815,L1816,L1817,L1818,L1819,L1820,L1821,L1822,L1823,L1824,L1825,L1826,L1827,L1828,L1829,L1830,L1831,L1832,L1833,L1834,L1835,L1836,L1837,L1838,L1839,L1840,L1841,L1842,L1843,L1844,L1845,L1846,L1847,L1848,L1849,L1850,L1851,L1852,L1853,L1854,L1855,L1856,L1857,L1858,L1859,L1860,L1861,L1862,L1863,L1864,L1865,L1866,L1867,L1868,L1869,L1870,L1871,L1872,L1873,L1874,L1875,L1876,L1877,L1878,L1879,L1880,L1881,L1882,L1883,L1884,L1885,L1886,L1887,L1888,L1889,L1890,L1891,L1892,L1893,L1894,L1895,L1896,L1897,L1898,L1899,L1900,L1901,L1902,L1903,L1904,L1905,L1906,L1907,L1908,L1909,L1910,L1911,L1912,L1913,L1914,L1915,L1916,L1917,L1918,L1919,L1920,L1921,L1922,L1923,L1924,L1925,L1926,L1927,L1928,L1929,L1930,L1931,L1932,L1933,L1934,L1935,L1936,L1937,L1938,L1939,L1940,L1941,L1942,L1943,L1944,L1945,L1946,L1947,L1948,L1949,L1950,L1951,L1952,L1953,L1954,L1955,L1956,L1957,L1958,L1959,L1960,L1961,L1962,L1963,L1964,L1965,L1966,L1967,L1968,L1969,L1970,L1971,L1972,L1973,L1974,L1975,L1976,L1977,L1978,L1979,L1980,L1981,L1982,L1983,L1984,L1985,L1986,L1987,L1988,L1989,L1990,L1991,L1992,L1993,L1994,L1995,L1996,L1997,L1998,L1999,L2000,L2001,L2002,L2003,L2004,L2005,L2006,L2007,L2008,L2009,L2010,L2011,L2012,L2013,L2014,L2015,L2016,L2017,L2018,L2019,L2020,L2021,L2022,L2023,L2024,L2025,L2026,L2027,L2028,L2029,L2030,L2031,L2032,L2033,L2034,L2035,L2036,L2037,L2038,L2039,L2040,L2041,L2042,L2043,L2044,L2045,L2046,L2047,L2048,L2049,L2050,L2051,L2052,L2053,L2054,L2055,L2056,L2057,L2058,L2059,L2060,L2061,L2062,L2063,L2064,L2065,L2066,L2067,L2068,L2069,L2070,L2071,L2072,L2073,L2074,L2075,L2076,L2077,L2078,L2079,L2080,L2081,L2082,L2083,L2084,L2085,L2086,L2087,L2088,L2089,L2090,L2091,L2092,L2093,L2094,L2095,L2096,L2097,L2098,L2099,L2100,L2101,L2102,L2103,L2104,L2105,L2106,L2107,L2108,L2109,L2110,L2111,L2112,L2113,L2114,L2115,L2116,L2117,L2118,L2119,L2120,L2121,L2122,L2123,L2124,L2125,L2126,L2127,L2128,L2129,L2130,L2131,L2132,L2133,L2134,L2135,L2136,L2137,L2138,L2139,L2140,L2141,L2142,L2143,L2144,L2145,L2146,L2147,L2148,L2149,L2150,L2151,L2152,L2153,L2154,L2155,L2156,L2157,L2158,L2159,L2160,L2161,L2162,L2163,L2164,L2165,L2166,L2167,L2168,L2169,L2170,L2171,L2172,L2173,L2174,L2175,L2176,L2177,L2178,L2179,L2180,L2181,L2182,L2183,L2184,L2185,L2186,L2187,L2188,L2189,L2190,L2191,L2192,L2193,L2194,L2195,L2196,L2197,L2198,L2199,L2200,L2201,L2202,L2203,L2204,L2205,L2206,L2207,L2208,L2209,L2210,L2211,L2212,L2213,L2214,L2215,L2216,L2217,L2218,L2219,L2220,L2221,L2222,L2223,L2224,L2225,L2226,L2227,L2228,L2229,L2230,L2231,L2232,L2233,L2234,L2235,L2236,L2237,L2238,L2239,L2240,L2241,L2242,L2243,L2244,L2245,L2246,L2247,L2248,L2249,L2250,L2251,L2252,L2253,L2254,L2255,L2256,L2257,L2258,L2259,L2260,L2261,L2262,L2263,L2264,L2265,L2266,L2267,L2268,L2269,L2270,L2271,L2272,L2273,L2274,L2275,L2276,L2277,L2278,L2279,L2280,L2281,L2282,L2283,L2284,L2285,L2286,L2287,L2288,L2289,L2290,L2291,L2292,L2293,L2294,L2295,L2296,L2297,L2298,L2299,L2300,L2301,L2302,L2303,L2304,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32,s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62,s63,s64,s65,s66,s67,s68,s69,s70,s71,s72,s73,s74,s75,s76,s77,s78,s79,s80,s81,s82,s83,s84,s85,s86,s87,s88,s89,s90,s91,s92,s93,s94,s95,s96,s97,s98,s99,s100,s101,s102,s103,s104,s105,s106,s107,s108,s109,s110,s111,s112,s113,s114,s115,s116,s117,s118,s119,s120,s121,s122,s123,s124,s125,s126,s127,s128,s129,s130,s131,s132,s133,s134,s135,s136,s137,s138,s139,s140,s141,s142,s143,s144,s145,s146,s147,s148,s149,s150,s151,s152,s153,s154,s155,s156,s157,s158,s159,s160,s161,s162,s163,s164,s165,s166,s167,s168,s169,s170,s171,s172,s173,s174,s175,s176,s177,s178,s179,s180,s181,s182,s183,s184,s185,s186,s187,s188,s189,s190,s191,s192,s193,s194,s195,s196,s197,s198,s199,s200,s201,s202,s203,s204,s205,s206,s207,s208,s209,s210,s211,s212,s213,s214,s215,s216,s217,s218,s219,s220,s221,s222,s223,s224,s225,s226,s227,s228,s229,s230,s231,s232,s233,s234,s235,s236,s237,s238,s239,s240,s241,s242,s243,s244,s245,s246,s247,s248,s249,s250,s251,s252,s253,s254,s255,s256,s257,s258,s259,s260,s261,s262,s263,s264,s265,s266,s267,s268,s269,s270,s271,s272,s273,s274,s275,s276,s277,s278,s279,s280,s281,s282,s283,s284,s285,s286,s287,s288,s289,s290,s291,s292,s293,s294,s295,s296,s297,s298,s299,s300,s301,s302,s303,s304,s305,s306,s307,s308,s309,s310,s311,s312,s313,s314,s315,s316,s317,s318,s319,s320,s321,s322,s323,s324,s325,s326,s327,s328,s329,s330,s331,s332,s333,s334,s335,s336,s337,s338,s339,s340,s341,s342,s343,s344,s345,s346,s347,s348,s349,s350,s351,s352,s353,s354,s355,s356,s357,s358,s359,s360,s361,s362,s363,s364,s365,s366,s367,s368,s369,s370,s371,s372,s373,s374,s375,s376,s377,s378,s379,s380,s381,s382,s383,s384,s385,s386,s387,s388,s389,s390,s391,s392,s393,s394,s395,s396,s397,s398,s399,s400,s401,s402,s403,s404,s405,s406,s407,s408,s409,s410,s411,s412,s413,s414,s415,s416,s417,s418,s419,s420,s421,s422,s423,s424,s425,s426,s427,s428,s429,s430,s431,s432,s433,s434,s435,s436,s437,s438,s439,s440,s441,s442,s443,s444,s445,s446,s447,s448,s449,s450,s451,s452,s453,s454,s455,s456,s457,s458,s459,s460,s461,s462,s463,s464,s465,s466,s467,s468,s469,s470,s471,s472,s473,s474,s475,s476,s477,s478,s479,s480,s481,s482,s483,s484,s485,s486,s487,s488,s489,s490,s491,s492,s493,s494,s495,s496,s497,s498,s499,s500,s501,s502,s503,s504,s505,s506,s507,s508,s509,s510,s511,s512,s513,s514,s515,s516,s517,s518,s519,s520,s521,s522,s523,s524,s525,s526,s527,s528,s529,s530,s531,s532,s533,s534,s535,s536,s537,s538,s539,s540,s541,s542,s543,s544,s545,s546,s547,s548,s549,s550,s551,s552,s553,s554,s555,s556,s557,s558,s559,s560,s561,s562,s563,s564,s565,s566,s567,s568,s569,s570,s571,s572,s573,s574,s575,s576,s577,s578,s579,s580,s581,s582,s583,s584,s585,s586,s587,s588,s589,s590,s591,s592,s593,s594,s595,s596,s597,s598,s599,s600,s601,s602,s603,s604,s605,s606,s607,s608,s609,s610,s611,s612,s613,s614,s615,s616,s617,s618,s619,s620,s621,s622,s623,s624,s625,s626,s627,s628,s629,s630,s631,s632,s633,s634,s635,s636,s637,s638,s639,s640,s641,s642,s643,s644,s645,s646,s647,s648,s649,s650,s651,s652,s653,s654,s655,s656,s657,s658,s659,s660,s661,s662,s663,s664,s665,s666,s667,s668,s669,s670,s671,s672,s673,s674,s675,s676,s677,s678,s679,s680,s681,s682,s683,s684,s685,s686,s687,s688,s689,s690,s691,s692,s693,s694,s695,s696,s697,s698,s699,s700,s701,s702,s703,s704,s705,s706,s707,s708,s709,s710,s711,s712,s713,s714,s715,s716,s717,s718,s719,s720,s721,s722,s723,s724,s725,s726,s727,s728,s729,s730,s731,s732,s733,s734,s735,s736,s737,s738,s739,s740,s741,s742,s743,s744,s745,s746,s747,s748,s749,s750,s751,s752,s753,s754,s755,s756,s757,s758,s759,s760,s761,s762,s763,s764,s765,s766,s767,s768,s769,s770,s771,s772,s773,s774,s775,s776,s777,s778,s779,s780,s781,s782,s783,s784,s785,s786,s787,s788,s789,s790,s791,s792,s793,s794,s795,s796,s797,s798,s799,s800,s801,s802,s803,s804,s805,s806,s807,s808,s809,s810,s811,s812,s813,s814,s815,s816,s817,s818,s819,s820,s821,s822,s823,s824,s825,s826,s827,s828,s829,s830,s831,s832,s833,s834,s835,s836,s837,s838,s839,s840,s841,s842,s843,s844,s845,s846,s847,s848,s849,s850,s851,s852,s853,s854,s855,s856,s857,s858,s859,s860,s861,s862,s863,s864,s865,s866,s867,s868,s869,s870,s871,s872,s873,s874,s875,s876,s877,s878,s879,s880,s881,s882,s883,s884,s885,s886,s887,s888,s889,s890,s891,s892,s893,s894,s895,s896,s897,s898,s899,s900,s901,s902,s903,s904,s905,s906,s907,s908,s909,s910,s911,s912,s913,s914,s915,s916,s917,s918,s919,s920,s921,s922,s923,s924,s925,s926,s927,s928,s929,s930,s931,s932,s933,s934,s935,s936,s937,s938,s939,s940,s941,s942,s943,s944,s945,s946,s947,s948,s949,s950,s951,s952,s953,s954,s955,s956,s957,s958,s959,s960,s961,s962,s963,s964,s965,s966,s967,s968,s969,s970,s971,s972,s973,s974,s975,s976,s977,s978,s979,s980,s981,s982,s983,s984,s985,s986,s987,s988,s989,s990,s991,s992,s993,s994,s995,s996,s997,s998,s999,s1000,s1001,s1002,s1003,s1004,s1005,s1006,s1007,s1008,s1009,s1010,s1011,s1012,s1013,s1014,s1015,s1016,s1017,s1018,s1019,s1020,s1021,s1022,s1023,s1024,s1025,s1026,s1027,s1028,s1029,s1030,s1031,s1032,s1033,s1034,s1035,s1036,s1037,s1038,s1039,s1040,s1041,s1042,s1043,s1044,s1045,s1046,s1047,s1048,s1049,s1050,s1051,s1052,s1053,s1054,s1055,s1056,s1057,s1058,s1059,s1060,s1061,s1062,s1063,s1064,s1065,s1066,s1067,s1068,s1069,s1070,s1071,s1072,s1073,s1074,s1075,s1076,s1077,s1078,s1079,s1080,s1081,s1082,s1083,s1084,s1085,s1086,s1087,s1088,s1089,s1090,s1091,s1092,s1093,s1094,s1095,s1096,s1097,s1098,s1099,s1100,s1101,s1102,s1103,s1104,s1105,s1106,s1107,s1108,s1109,s1110,s1111,s1112,s1113,s1114,s1115,s1116,s1117,s1118,s1119,s1120,s1121,s1122,s1123,s1124,s1125,s1126,s1127,s1128,s1129,s1130,s1131,s1132,s1133,s1134,s1135,s1136,s1137,s1138,s1139,s1140,s1141,s1142,s1143,s1144,s1145,s1146,s1147,s1148,s1149,s1150,s1151,s1152,s1153,s1154,s1155,s1156,s1157,s1158,s1159,s1160,s1161,s1162,s1163,s1164,s1165,s1166,s1167,s1168,s1169,s1170,s1171,s1172,s1173,s1174,s1175,s1176,s1177,s1178,s1179,s1180,s1181,s1182,s1183,s1184,s1185,s1186,s1187,s1188,s1189,s1190,s1191,s1192,s1193,s1194,s1195,s1196,s1197,s1198,s1199,s1200,s1201,s1202,s1203,s1204,s1205,s1206,s1207,s1208,s1209,s1210,s1211,s1212,s1213,s1214,s1215,s1216,s1217,s1218,s1219,s1220,s1221,s1222,s1223,s1224,s1225,s1226,s1227,s1228,s1229,s1230,s1231,s1232,s1233,s1234,s1235,s1236,s1237,s1238,s1239,s1240,s1241,s1242,s1243,s1244,s1245,s1246,s1247,s1248,s1249,s1250,s1251,s1252,s1253,s1254,s1255,s1256,s1257,s1258,s1259,s1260,s1261,s1262,s1263,s1264,s1265,s1266,s1267,s1268,s1269,s1270,s1271,s1272,s1273,s1274,s1275,s1276,s1277,s1278,s1279,s1280,s1281,s1282,s1283,s1284,s1285,s1286,s1287,s1288,s1289,s1290,s1291,s1292,s1293,s1294,s1295,s1296,s1297,s1298,s1299,s1300,s1301,s1302,s1303,s1304,s1305,s1306,s1307,s1308,s1309,s1310,s1311,s1312,s1313,s1314,s1315,s1316,s1317,s1318,s1319,s1320,s1321,s1322,s1323,s1324,s1325,s1326,s1327,s1328,s1329,s1330,s1331,s1332,s1333,s1334,s1335,s1336,s1337,s1338,s1339,s1340,s1341,s1342,s1343,s1344,s1345,s1346,s1347,s1348,s1349,s1350,s1351,s1352,s1353,s1354,s1355,s1356,s1357,s1358,s1359,s1360,s1361,s1362,s1363,s1364,s1365,s1366,s1367,s1368,s1369,s1370,s1371,s1372,s1373,s1374,s1375,s1376,s1377,s1378,s1379,s1380,s1381,s1382,s1383,s1384,s1385,s1386,s1387,s1388,s1389,s1390,s1391,s1392,s1393,s1394,s1395,s1396,s1397,s1398,s1399,s1400,s1401,s1402,s1403,s1404,s1405,s1406,s1407,s1408,s1409,s1410,s1411,s1412,s1413,s1414,s1415,s1416,s1417,s1418,s1419,s1420,s1421,s1422,s1423,s1424,s1425,s1426,s1427,s1428,s1429,s1430,s1431,s1432,s1433,s1434,s1435,s1436,s1437,s1438,s1439,s1440,s1441,s1442,s1443,s1444,s1445,s1446,s1447,s1448,s1449,s1450,s1451,s1452,s1453,s1454,s1455,s1456,s1457,s1458,s1459,s1460,s1461,s1462,s1463,s1464,s1465,s1466,s1467,s1468,s1469,s1470,s1471,s1472,s1473,s1474,s1475,s1476,s1477,s1478,s1479,s1480,s1481,s1482,s1483,s1484,s1485,s1486,s1487,s1488,s1489,s1490,s1491,s1492,s1493,s1494,s1495,s1496,s1497,s1498,s1499,s1500,s1501,s1502,s1503,s1504,s1505,s1506,s1507,s1508,s1509,s1510,s1511,s1512,s1513,s1514,s1515,s1516,s1517,s1518,s1519,s1520,s1521,s1522,s1523,s1524,s1525,s1526,s1527,s1528,s1529,s1530,s1531,s1532,s1533,s1534,s1535,s1536,s1537,s1538,s1539,s1540,s1541,s1542,s1543,s1544,s1545,s1546,s1547,s1548,s1549,s1550,s1551,s1552,s1553,s1554,s1555,s1556,s1557,s1558,s1559,s1560,s1561,s1562,s1563,s1564,s1565,s1566,s1567,s1568,s1569,s1570,s1571,s1572,s1573,s1574,s1575,s1576,s1577,s1578,s1579,s1580,s1581,s1582,s1583,s1584,s1585,s1586,s1587,s1588,s1589,s1590,s1591,s1592,s1593,s1594,s1595,s1596,s1597,s1598,s1599,s1600,s1601,s1602,s1603,s1604,s1605,s1606,s1607,s1608,s1609,s1610,s1611,s1612,s1613,s1614,s1615,s1616,s1617,s1618,s1619,s1620,s1621,s1622,s1623,s1624,s1625,s1626,s1627,s1628,s1629,s1630,s1631,s1632,s1633,s1634,s1635,s1636,s1637,s1638,s1639,s1640,s1641,s1642,s1643,s1644,s1645,s1646,s1647,s1648,s1649,s1650,s1651,s1652,s1653,s1654,s1655,s1656,s1657,s1658,s1659,s1660,s1661,s1662,s1663,s1664,s1665,s1666,s1667,s1668,s1669,s1670,s1671,s1672,s1673,s1674,s1675,s1676,s1677,s1678,s1679,s1680,s1681,s1682,s1683,s1684,s1685,s1686,s1687,s1688,s1689,s1690,s1691,s1692,s1693,s1694,s1695,s1696,s1697,s1698,s1699,s1700,s1701,s1702,s1703,s1704,s1705,s1706,s1707,s1708,s1709,s1710,s1711,s1712,s1713,s1714,s1715,s1716,s1717,s1718,s1719,s1720,s1721,s1722,s1723,s1724,s1725,s1726,s1727,s1728,s1729,s1730,s1731,s1732,s1733,s1734,s1735,s1736,s1737,s1738,s1739,s1740,s1741,s1742,s1743,s1744,s1745,s1746,s1747,s1748,s1749,s1750,s1751,s1752,s1753,s1754,s1755,s1756,s1757,s1758,s1759,s1760,s1761,s1762,s1763,s1764,s1765,s1766,s1767,s1768,s1769,s1770,s1771,s1772,s1773,s1774,s1775,s1776,s1777,s1778,s1779,s1780,s1781,s1782,s1783,s1784,s1785,s1786,s1787,s1788,s1789,s1790,s1791,s1792,s1793,s1794,s1795,s1796,s1797,s1798,s1799,s1800,s1801,s1802,s1803,s1804,s1805,s1806,s1807,s1808,s1809,s1810,s1811,s1812,s1813,s1814,s1815,s1816,s1817,s1818,s1819,s1820,s1821,s1822,s1823,s1824,s1825,s1826,s1827,s1828,s1829,s1830,s1831,s1832,s1833,s1834,s1835,s1836,s1837,s1838,s1839,s1840,s1841,s1842,s1843,s1844,s1845,s1846,s1847,s1848,s1849,s1850,s1851,s1852,s1853,s1854,s1855,s1856,s1857,s1858,s1859,s1860,s1861,s1862,s1863,s1864,s1865,s1866,s1867,s1868,s1869,s1870,s1871,s1872,s1873,s1874,s1875,s1876,s1877,s1878,s1879,s1880,s1881,s1882,s1883,s1884,s1885,s1886,s1887,s1888,s1889,s1890,s1891,s1892,s1893,s1894,s1895,s1896,s1897,s1898,s1899,s1900,s1901,s1902,s1903,s1904,s1905,s1906,s1907,s1908,s1909,s1910,s1911,s1912,s1913,s1914,s1915,s1916,s1917,s1918,s1919,s1920,s1921,s1922,s1923,s1924,s1925,s1926,s1927,s1928,s1929,s1930,s1931,s1932,s1933,s1934,s1935,s1936,s1937,s1938,s1939,s1940,s1941,s1942,s1943,s1944,s1945,s1946,s1947,s1948,s1949,s1950,s1951,s1952,s1953,s1954,s1955,s1956,s1957,s1958,s1959,s1960,s1961,s1962,s1963,s1964,s1965,s1966,s1967,s1968,s1969,s1970,s1971,s1972,s1973,s1974,s1975,s1976,s1977,s1978,s1979,s1980,s1981,s1982,s1983,s1984,s1985,s1986,s1987,s1988,s1989,s1990,s1991,s1992,s1993,s1994,s1995,s1996,s1997,s1998,s1999,s2000,s2001,s2002,s2003,s2004,s2005,s2006,s2007,s2008,s2009,s2010,s2011,s2012,s2013,s2014,s2015,s2016,s2017,s2018,s2019,s2020,s2021,s2022,s2023,s2024,s2025,s2026,s2027,s2028,s2029,s2030,s2031,s2032,s2033,s2034,s2035,s2036,s2037,s2038,s2039,s2040,s2041,s2042,s2043,s2044,s2045,s2046,s2047,s2048,s2049,s2050,s2051,s2052,s2053,s2054,s2055,s2056,s2057,s2058,s2059,s2060,s2061,s2062,s2063,s2064,s2065,s2066,s2067,s2068,s2069,s2070,s2071,s2072,s2073,s2074,s2075,s2076,s2077,s2078,s2079,s2080,s2081,s2082,s2083,s2084,s2085,s2086,s2087,s2088,s2089,s2090,s2091,s2092,s2093,s2094,s2095,s2096,s2097,s2098,s2099,s2100,s2101,s2102,s2103,s2104,s2105,s2106,s2107,s2108,s2109,s2110,s2111,s2112,s2113,s2114,s2115,s2116,s2117,s2118,s2119,s2120,s2121,s2122,s2123,s2124,s2125,s2126,s2127,s2128,s2129,s2130,s2131,s2132,s2133,s2134,s2135,s2136,s2137,s2138,s2139,s2140,s2141,s2142,s2143,s2144,s2145,s2146,s2147,s2148,s2149,s2150,s2151,s2152,s2153,s2154,s2155,s2156,s2157,s2158,s2159,s2160,s2161,s2162,s2163,s2164,s2165,s2166,s2167,s2168,s2169,s2170,s2171,s2172,s2173,s2174,s2175,s2176,s2177,s2178,s2179,s2180,s2181,s2182,s2183,s2184,s2185,s2186,s2187,s2188,s2189,s2190,s2191,s2192,s2193,s2194,s2195,s2196,s2197,s2198,s2199,s2200,s2201,s2202,s2203,s2204,s2205,s2206,s2207,s2208,s2209,s2210,s2211,s2212,s2213,s2214,s2215,s2216,s2217,s2218,s2219,s2220,s2221,s2222,s2223,s2224,s2225,s2226,s2227,s2228,s2229,s2230,s2231,s2232,s2233,s2234,s2235,s2236,s2237,s2238,s2239,s2240,s2241,s2242,s2243,s2244,s2245,s2246,s2247,s2248,s2249,s2250,s2251,s2252,s2253,s2254,s2255,s2256,s2257,s2258,s2259,s2260,s2261,s2262,s2263,s2264,s2265,s2266,s2267,s2268,s2269,s2270,s2271,s2272,s2273,s2274,s2275,s2276,s2277,s2278,s2279,s2280,s2281,s2282,s2283,s2284,s2285,s2286,s2287,s2288,s2289,s2290,s2291,s2292,s2293,s2294,s2295,s2296,s2297,s2298,s2299,s2300,s2301,s2302,s2303,s2304,x_x,y_y);

Z1<=s1;
Z2<=s2;
Z3<=s3;
Z4<=s4;
Z5<=s5;
Z6<=s6;
Z7<=s7;
Z8<=s8;
Z9<=s9;
Z10<=s10;
Z11<=s11;
Z12<=s12;
Z13<=s13;
Z14<=s14;
Z15<=s15;
Z16<=s16;
Z17<=s17;
Z18<=s18;
Z19<=s19;
Z20<=s20;
Z21<=s21;
Z22<=s22;
Z23<=s23;
Z24<=s24;
Z25<=s25;
Z26<=s26;
Z27<=s27;
Z28<=s28;
Z29<=s29;
Z30<=s30;
Z31<=s31;
Z32<=s32;
Z33<=s33;
Z34<=s34;
Z35<=s35;
Z36<=s36;
Z37<=s37;
Z38<=s38;
Z39<=s39;
Z40<=s40;
Z41<=s41;
Z42<=s42;
Z43<=s43;
Z44<=s44;
Z45<=s45;
Z46<=s46;
Z47<=s47;
Z48<=s48;
Z49<=s49;
Z50<=s50;
Z51<=s51;
Z52<=s52;
Z53<=s53;
Z54<=s54;
Z55<=s55;
Z56<=s56;
Z57<=s57;
Z58<=s58;
Z59<=s59;
Z60<=s60;
Z61<=s61;
Z62<=s62;
Z63<=s63;
Z64<=s64;
Z65<=s65;
Z66<=s66;
Z67<=s67;
Z68<=s68;
Z69<=s69;
Z70<=s70;
Z71<=s71;
Z72<=s72;
Z73<=s73;
Z74<=s74;
Z75<=s75;
Z76<=s76;
Z77<=s77;
Z78<=s78;
Z79<=s79;
Z80<=s80;
Z81<=s81;
Z82<=s82;
Z83<=s83;
Z84<=s84;
Z85<=s85;
Z86<=s86;
Z87<=s87;
Z88<=s88;
Z89<=s89;
Z90<=s90;
Z91<=s91;
Z92<=s92;
Z93<=s93;
Z94<=s94;
Z95<=s95;
Z96<=s96;
Z97<=s97;
Z98<=s98;
Z99<=s99;
Z100<=s100;
Z101<=s101;
Z102<=s102;
Z103<=s103;
Z104<=s104;
Z105<=s105;
Z106<=s106;
Z107<=s107;
Z108<=s108;
Z109<=s109;
Z110<=s110;
Z111<=s111;
Z112<=s112;
Z113<=s113;
Z114<=s114;
Z115<=s115;
Z116<=s116;
Z117<=s117;
Z118<=s118;
Z119<=s119;
Z120<=s120;
Z121<=s121;
Z122<=s122;
Z123<=s123;
Z124<=s124;
Z125<=s125;
Z126<=s126;
Z127<=s127;
Z128<=s128;
Z129<=s129;
Z130<=s130;
Z131<=s131;
Z132<=s132;
Z133<=s133;
Z134<=s134;
Z135<=s135;
Z136<=s136;
Z137<=s137;
Z138<=s138;
Z139<=s139;
Z140<=s140;
Z141<=s141;
Z142<=s142;
Z143<=s143;
Z144<=s144;
Z145<=s145;
Z146<=s146;
Z147<=s147;
Z148<=s148;
Z149<=s149;
Z150<=s150;
Z151<=s151;
Z152<=s152;
Z153<=s153;
Z154<=s154;
Z155<=s155;
Z156<=s156;
Z157<=s157;
Z158<=s158;
Z159<=s159;
Z160<=s160;
Z161<=s161;
Z162<=s162;
Z163<=s163;
Z164<=s164;
Z165<=s165;
Z166<=s166;
Z167<=s167;
Z168<=s168;
Z169<=s169;
Z170<=s170;
Z171<=s171;
Z172<=s172;
Z173<=s173;
Z174<=s174;
Z175<=s175;
Z176<=s176;
Z177<=s177;
Z178<=s178;
Z179<=s179;
Z180<=s180;
Z181<=s181;
Z182<=s182;
Z183<=s183;
Z184<=s184;
Z185<=s185;
Z186<=s186;
Z187<=s187;
Z188<=s188;
Z189<=s189;
Z190<=s190;
Z191<=s191;
Z192<=s192;
Z193<=s193;
Z194<=s194;
Z195<=s195;
Z196<=s196;
Z197<=s197;
Z198<=s198;
Z199<=s199;
Z200<=s200;
Z201<=s201;
Z202<=s202;
Z203<=s203;
Z204<=s204;
Z205<=s205;
Z206<=s206;
Z207<=s207;
Z208<=s208;
Z209<=s209;
Z210<=s210;
Z211<=s211;
Z212<=s212;
Z213<=s213;
Z214<=s214;
Z215<=s215;
Z216<=s216;
Z217<=s217;
Z218<=s218;
Z219<=s219;
Z220<=s220;
Z221<=s221;
Z222<=s222;
Z223<=s223;
Z224<=s224;
Z225<=s225;
Z226<=s226;
Z227<=s227;
Z228<=s228;
Z229<=s229;
Z230<=s230;
Z231<=s231;
Z232<=s232;
Z233<=s233;
Z234<=s234;
Z235<=s235;
Z236<=s236;
Z237<=s237;
Z238<=s238;
Z239<=s239;
Z240<=s240;
Z241<=s241;
Z242<=s242;
Z243<=s243;
Z244<=s244;
Z245<=s245;
Z246<=s246;
Z247<=s247;
Z248<=s248;
Z249<=s249;
Z250<=s250;
Z251<=s251;
Z252<=s252;
Z253<=s253;
Z254<=s254;
Z255<=s255;
Z256<=s256;
Z257<=s257;
Z258<=s258;
Z259<=s259;
Z260<=s260;
Z261<=s261;
Z262<=s262;
Z263<=s263;
Z264<=s264;
Z265<=s265;
Z266<=s266;
Z267<=s267;
Z268<=s268;
Z269<=s269;
Z270<=s270;
Z271<=s271;
Z272<=s272;
Z273<=s273;
Z274<=s274;
Z275<=s275;
Z276<=s276;
Z277<=s277;
Z278<=s278;
Z279<=s279;
Z280<=s280;
Z281<=s281;
Z282<=s282;
Z283<=s283;
Z284<=s284;
Z285<=s285;
Z286<=s286;
Z287<=s287;
Z288<=s288;
Z289<=s289;
Z290<=s290;
Z291<=s291;
Z292<=s292;
Z293<=s293;
Z294<=s294;
Z295<=s295;
Z296<=s296;
Z297<=s297;
Z298<=s298;
Z299<=s299;
Z300<=s300;
Z301<=s301;
Z302<=s302;
Z303<=s303;
Z304<=s304;
Z305<=s305;
Z306<=s306;
Z307<=s307;
Z308<=s308;
Z309<=s309;
Z310<=s310;
Z311<=s311;
Z312<=s312;
Z313<=s313;
Z314<=s314;
Z315<=s315;
Z316<=s316;
Z317<=s317;
Z318<=s318;
Z319<=s319;
Z320<=s320;
Z321<=s321;
Z322<=s322;
Z323<=s323;
Z324<=s324;
Z325<=s325;
Z326<=s326;
Z327<=s327;
Z328<=s328;
Z329<=s329;
Z330<=s330;
Z331<=s331;
Z332<=s332;
Z333<=s333;
Z334<=s334;
Z335<=s335;
Z336<=s336;
Z337<=s337;
Z338<=s338;
Z339<=s339;
Z340<=s340;
Z341<=s341;
Z342<=s342;
Z343<=s343;
Z344<=s344;
Z345<=s345;
Z346<=s346;
Z347<=s347;
Z348<=s348;
Z349<=s349;
Z350<=s350;
Z351<=s351;
Z352<=s352;
Z353<=s353;
Z354<=s354;
Z355<=s355;
Z356<=s356;
Z357<=s357;
Z358<=s358;
Z359<=s359;
Z360<=s360;
Z361<=s361;
Z362<=s362;
Z363<=s363;
Z364<=s364;
Z365<=s365;
Z366<=s366;
Z367<=s367;
Z368<=s368;
Z369<=s369;
Z370<=s370;
Z371<=s371;
Z372<=s372;
Z373<=s373;
Z374<=s374;
Z375<=s375;
Z376<=s376;
Z377<=s377;
Z378<=s378;
Z379<=s379;
Z380<=s380;
Z381<=s381;
Z382<=s382;
Z383<=s383;
Z384<=s384;
Z385<=s385;
Z386<=s386;
Z387<=s387;
Z388<=s388;
Z389<=s389;
Z390<=s390;
Z391<=s391;
Z392<=s392;
Z393<=s393;
Z394<=s394;
Z395<=s395;
Z396<=s396;
Z397<=s397;
Z398<=s398;
Z399<=s399;
Z400<=s400;
Z401<=s401;
Z402<=s402;
Z403<=s403;
Z404<=s404;
Z405<=s405;
Z406<=s406;
Z407<=s407;
Z408<=s408;
Z409<=s409;
Z410<=s410;
Z411<=s411;
Z412<=s412;
Z413<=s413;
Z414<=s414;
Z415<=s415;
Z416<=s416;
Z417<=s417;
Z418<=s418;
Z419<=s419;
Z420<=s420;
Z421<=s421;
Z422<=s422;
Z423<=s423;
Z424<=s424;
Z425<=s425;
Z426<=s426;
Z427<=s427;
Z428<=s428;
Z429<=s429;
Z430<=s430;
Z431<=s431;
Z432<=s432;
Z433<=s433;
Z434<=s434;
Z435<=s435;
Z436<=s436;
Z437<=s437;
Z438<=s438;
Z439<=s439;
Z440<=s440;
Z441<=s441;
Z442<=s442;
Z443<=s443;
Z444<=s444;
Z445<=s445;
Z446<=s446;
Z447<=s447;
Z448<=s448;
Z449<=s449;
Z450<=s450;
Z451<=s451;
Z452<=s452;
Z453<=s453;
Z454<=s454;
Z455<=s455;
Z456<=s456;
Z457<=s457;
Z458<=s458;
Z459<=s459;
Z460<=s460;
Z461<=s461;
Z462<=s462;
Z463<=s463;
Z464<=s464;
Z465<=s465;
Z466<=s466;
Z467<=s467;
Z468<=s468;
Z469<=s469;
Z470<=s470;
Z471<=s471;
Z472<=s472;
Z473<=s473;
Z474<=s474;
Z475<=s475;
Z476<=s476;
Z477<=s477;
Z478<=s478;
Z479<=s479;
Z480<=s480;
Z481<=s481;
Z482<=s482;
Z483<=s483;
Z484<=s484;
Z485<=s485;
Z486<=s486;
Z487<=s487;
Z488<=s488;
Z489<=s489;
Z490<=s490;
Z491<=s491;
Z492<=s492;
Z493<=s493;
Z494<=s494;
Z495<=s495;
Z496<=s496;
Z497<=s497;
Z498<=s498;
Z499<=s499;
Z500<=s500;
Z501<=s501;
Z502<=s502;
Z503<=s503;
Z504<=s504;
Z505<=s505;
Z506<=s506;
Z507<=s507;
Z508<=s508;
Z509<=s509;
Z510<=s510;
Z511<=s511;
Z512<=s512;
Z513<=s513;
Z514<=s514;
Z515<=s515;
Z516<=s516;
Z517<=s517;
Z518<=s518;
Z519<=s519;
Z520<=s520;
Z521<=s521;
Z522<=s522;
Z523<=s523;
Z524<=s524;
Z525<=s525;
Z526<=s526;
Z527<=s527;
Z528<=s528;
Z529<=s529;
Z530<=s530;
Z531<=s531;
Z532<=s532;
Z533<=s533;
Z534<=s534;
Z535<=s535;
Z536<=s536;
Z537<=s537;
Z538<=s538;
Z539<=s539;
Z540<=s540;
Z541<=s541;
Z542<=s542;
Z543<=s543;
Z544<=s544;
Z545<=s545;
Z546<=s546;
Z547<=s547;
Z548<=s548;
Z549<=s549;
Z550<=s550;
Z551<=s551;
Z552<=s552;
Z553<=s553;
Z554<=s554;
Z555<=s555;
Z556<=s556;
Z557<=s557;
Z558<=s558;
Z559<=s559;
Z560<=s560;
Z561<=s561;
Z562<=s562;
Z563<=s563;
Z564<=s564;
Z565<=s565;
Z566<=s566;
Z567<=s567;
Z568<=s568;
Z569<=s569;
Z570<=s570;
Z571<=s571;
Z572<=s572;
Z573<=s573;
Z574<=s574;
Z575<=s575;
Z576<=s576;
Z577<=s577;
Z578<=s578;
Z579<=s579;
Z580<=s580;
Z581<=s581;
Z582<=s582;
Z583<=s583;
Z584<=s584;
Z585<=s585;
Z586<=s586;
Z587<=s587;
Z588<=s588;
Z589<=s589;
Z590<=s590;
Z591<=s591;
Z592<=s592;
Z593<=s593;
Z594<=s594;
Z595<=s595;
Z596<=s596;
Z597<=s597;
Z598<=s598;
Z599<=s599;
Z600<=s600;
Z601<=s601;
Z602<=s602;
Z603<=s603;
Z604<=s604;
Z605<=s605;
Z606<=s606;
Z607<=s607;
Z608<=s608;
Z609<=s609;
Z610<=s610;
Z611<=s611;
Z612<=s612;
Z613<=s613;
Z614<=s614;
Z615<=s615;
Z616<=s616;
Z617<=s617;
Z618<=s618;
Z619<=s619;
Z620<=s620;
Z621<=s621;
Z622<=s622;
Z623<=s623;
Z624<=s624;
Z625<=s625;
Z626<=s626;
Z627<=s627;
Z628<=s628;
Z629<=s629;
Z630<=s630;
Z631<=s631;
Z632<=s632;
Z633<=s633;
Z634<=s634;
Z635<=s635;
Z636<=s636;
Z637<=s637;
Z638<=s638;
Z639<=s639;
Z640<=s640;
Z641<=s641;
Z642<=s642;
Z643<=s643;
Z644<=s644;
Z645<=s645;
Z646<=s646;
Z647<=s647;
Z648<=s648;
Z649<=s649;
Z650<=s650;
Z651<=s651;
Z652<=s652;
Z653<=s653;
Z654<=s654;
Z655<=s655;
Z656<=s656;
Z657<=s657;
Z658<=s658;
Z659<=s659;
Z660<=s660;
Z661<=s661;
Z662<=s662;
Z663<=s663;
Z664<=s664;
Z665<=s665;
Z666<=s666;
Z667<=s667;
Z668<=s668;
Z669<=s669;
Z670<=s670;
Z671<=s671;
Z672<=s672;
Z673<=s673;
Z674<=s674;
Z675<=s675;
Z676<=s676;
Z677<=s677;
Z678<=s678;
Z679<=s679;
Z680<=s680;
Z681<=s681;
Z682<=s682;
Z683<=s683;
Z684<=s684;
Z685<=s685;
Z686<=s686;
Z687<=s687;
Z688<=s688;
Z689<=s689;
Z690<=s690;
Z691<=s691;
Z692<=s692;
Z693<=s693;
Z694<=s694;
Z695<=s695;
Z696<=s696;
Z697<=s697;
Z698<=s698;
Z699<=s699;
Z700<=s700;
Z701<=s701;
Z702<=s702;
Z703<=s703;
Z704<=s704;
Z705<=s705;
Z706<=s706;
Z707<=s707;
Z708<=s708;
Z709<=s709;
Z710<=s710;
Z711<=s711;
Z712<=s712;
Z713<=s713;
Z714<=s714;
Z715<=s715;
Z716<=s716;
Z717<=s717;
Z718<=s718;
Z719<=s719;
Z720<=s720;
Z721<=s721;
Z722<=s722;
Z723<=s723;
Z724<=s724;
Z725<=s725;
Z726<=s726;
Z727<=s727;
Z728<=s728;
Z729<=s729;
Z730<=s730;
Z731<=s731;
Z732<=s732;
Z733<=s733;
Z734<=s734;
Z735<=s735;
Z736<=s736;
Z737<=s737;
Z738<=s738;
Z739<=s739;
Z740<=s740;
Z741<=s741;
Z742<=s742;
Z743<=s743;
Z744<=s744;
Z745<=s745;
Z746<=s746;
Z747<=s747;
Z748<=s748;
Z749<=s749;
Z750<=s750;
Z751<=s751;
Z752<=s752;
Z753<=s753;
Z754<=s754;
Z755<=s755;
Z756<=s756;
Z757<=s757;
Z758<=s758;
Z759<=s759;
Z760<=s760;
Z761<=s761;
Z762<=s762;
Z763<=s763;
Z764<=s764;
Z765<=s765;
Z766<=s766;
Z767<=s767;
Z768<=s768;
Z769<=s769;
Z770<=s770;
Z771<=s771;
Z772<=s772;
Z773<=s773;
Z774<=s774;
Z775<=s775;
Z776<=s776;
Z777<=s777;
Z778<=s778;
Z779<=s779;
Z780<=s780;
Z781<=s781;
Z782<=s782;
Z783<=s783;
Z784<=s784;
Z785<=s785;
Z786<=s786;
Z787<=s787;
Z788<=s788;
Z789<=s789;
Z790<=s790;
Z791<=s791;
Z792<=s792;
Z793<=s793;
Z794<=s794;
Z795<=s795;
Z796<=s796;
Z797<=s797;
Z798<=s798;
Z799<=s799;
Z800<=s800;
Z801<=s801;
Z802<=s802;
Z803<=s803;
Z804<=s804;
Z805<=s805;
Z806<=s806;
Z807<=s807;
Z808<=s808;
Z809<=s809;
Z810<=s810;
Z811<=s811;
Z812<=s812;
Z813<=s813;
Z814<=s814;
Z815<=s815;
Z816<=s816;
Z817<=s817;
Z818<=s818;
Z819<=s819;
Z820<=s820;
Z821<=s821;
Z822<=s822;
Z823<=s823;
Z824<=s824;
Z825<=s825;
Z826<=s826;
Z827<=s827;
Z828<=s828;
Z829<=s829;
Z830<=s830;
Z831<=s831;
Z832<=s832;
Z833<=s833;
Z834<=s834;
Z835<=s835;
Z836<=s836;
Z837<=s837;
Z838<=s838;
Z839<=s839;
Z840<=s840;
Z841<=s841;
Z842<=s842;
Z843<=s843;
Z844<=s844;
Z845<=s845;
Z846<=s846;
Z847<=s847;
Z848<=s848;
Z849<=s849;
Z850<=s850;
Z851<=s851;
Z852<=s852;
Z853<=s853;
Z854<=s854;
Z855<=s855;
Z856<=s856;
Z857<=s857;
Z858<=s858;
Z859<=s859;
Z860<=s860;
Z861<=s861;
Z862<=s862;
Z863<=s863;
Z864<=s864;
Z865<=s865;
Z866<=s866;
Z867<=s867;
Z868<=s868;
Z869<=s869;
Z870<=s870;
Z871<=s871;
Z872<=s872;
Z873<=s873;
Z874<=s874;
Z875<=s875;
Z876<=s876;
Z877<=s877;
Z878<=s878;
Z879<=s879;
Z880<=s880;
Z881<=s881;
Z882<=s882;
Z883<=s883;
Z884<=s884;
Z885<=s885;
Z886<=s886;
Z887<=s887;
Z888<=s888;
Z889<=s889;
Z890<=s890;
Z891<=s891;
Z892<=s892;
Z893<=s893;
Z894<=s894;
Z895<=s895;
Z896<=s896;
Z897<=s897;
Z898<=s898;
Z899<=s899;
Z900<=s900;
Z901<=s901;
Z902<=s902;
Z903<=s903;
Z904<=s904;
Z905<=s905;
Z906<=s906;
Z907<=s907;
Z908<=s908;
Z909<=s909;
Z910<=s910;
Z911<=s911;
Z912<=s912;
Z913<=s913;
Z914<=s914;
Z915<=s915;
Z916<=s916;
Z917<=s917;
Z918<=s918;
Z919<=s919;
Z920<=s920;
Z921<=s921;
Z922<=s922;
Z923<=s923;
Z924<=s924;
Z925<=s925;
Z926<=s926;
Z927<=s927;
Z928<=s928;
Z929<=s929;
Z930<=s930;
Z931<=s931;
Z932<=s932;
Z933<=s933;
Z934<=s934;
Z935<=s935;
Z936<=s936;
Z937<=s937;
Z938<=s938;
Z939<=s939;
Z940<=s940;
Z941<=s941;
Z942<=s942;
Z943<=s943;
Z944<=s944;
Z945<=s945;
Z946<=s946;
Z947<=s947;
Z948<=s948;
Z949<=s949;
Z950<=s950;
Z951<=s951;
Z952<=s952;
Z953<=s953;
Z954<=s954;
Z955<=s955;
Z956<=s956;
Z957<=s957;
Z958<=s958;
Z959<=s959;
Z960<=s960;
Z961<=s961;
Z962<=s962;
Z963<=s963;
Z964<=s964;
Z965<=s965;
Z966<=s966;
Z967<=s967;
Z968<=s968;
Z969<=s969;
Z970<=s970;
Z971<=s971;
Z972<=s972;
Z973<=s973;
Z974<=s974;
Z975<=s975;
Z976<=s976;
Z977<=s977;
Z978<=s978;
Z979<=s979;
Z980<=s980;
Z981<=s981;
Z982<=s982;
Z983<=s983;
Z984<=s984;
Z985<=s985;
Z986<=s986;
Z987<=s987;
Z988<=s988;
Z989<=s989;
Z990<=s990;
Z991<=s991;
Z992<=s992;
Z993<=s993;
Z994<=s994;
Z995<=s995;
Z996<=s996;
Z997<=s997;
Z998<=s998;
Z999<=s999;
Z1000<=s1000;
Z1001<=s1001;
Z1002<=s1002;
Z1003<=s1003;
Z1004<=s1004;
Z1005<=s1005;
Z1006<=s1006;
Z1007<=s1007;
Z1008<=s1008;
Z1009<=s1009;
Z1010<=s1010;
Z1011<=s1011;
Z1012<=s1012;
Z1013<=s1013;
Z1014<=s1014;
Z1015<=s1015;
Z1016<=s1016;
Z1017<=s1017;
Z1018<=s1018;
Z1019<=s1019;
Z1020<=s1020;
Z1021<=s1021;
Z1022<=s1022;
Z1023<=s1023;
Z1024<=s1024;
Z1025<=s1025;
Z1026<=s1026;
Z1027<=s1027;
Z1028<=s1028;
Z1029<=s1029;
Z1030<=s1030;
Z1031<=s1031;
Z1032<=s1032;
Z1033<=s1033;
Z1034<=s1034;
Z1035<=s1035;
Z1036<=s1036;
Z1037<=s1037;
Z1038<=s1038;
Z1039<=s1039;
Z1040<=s1040;
Z1041<=s1041;
Z1042<=s1042;
Z1043<=s1043;
Z1044<=s1044;
Z1045<=s1045;
Z1046<=s1046;
Z1047<=s1047;
Z1048<=s1048;
Z1049<=s1049;
Z1050<=s1050;
Z1051<=s1051;
Z1052<=s1052;
Z1053<=s1053;
Z1054<=s1054;
Z1055<=s1055;
Z1056<=s1056;
Z1057<=s1057;
Z1058<=s1058;
Z1059<=s1059;
Z1060<=s1060;
Z1061<=s1061;
Z1062<=s1062;
Z1063<=s1063;
Z1064<=s1064;
Z1065<=s1065;
Z1066<=s1066;
Z1067<=s1067;
Z1068<=s1068;
Z1069<=s1069;
Z1070<=s1070;
Z1071<=s1071;
Z1072<=s1072;
Z1073<=s1073;
Z1074<=s1074;
Z1075<=s1075;
Z1076<=s1076;
Z1077<=s1077;
Z1078<=s1078;
Z1079<=s1079;
Z1080<=s1080;
Z1081<=s1081;
Z1082<=s1082;
Z1083<=s1083;
Z1084<=s1084;
Z1085<=s1085;
Z1086<=s1086;
Z1087<=s1087;
Z1088<=s1088;
Z1089<=s1089;
Z1090<=s1090;
Z1091<=s1091;
Z1092<=s1092;
Z1093<=s1093;
Z1094<=s1094;
Z1095<=s1095;
Z1096<=s1096;
Z1097<=s1097;
Z1098<=s1098;
Z1099<=s1099;
Z1100<=s1100;
Z1101<=s1101;
Z1102<=s1102;
Z1103<=s1103;
Z1104<=s1104;
Z1105<=s1105;
Z1106<=s1106;
Z1107<=s1107;
Z1108<=s1108;
Z1109<=s1109;
Z1110<=s1110;
Z1111<=s1111;
Z1112<=s1112;
Z1113<=s1113;
Z1114<=s1114;
Z1115<=s1115;
Z1116<=s1116;
Z1117<=s1117;
Z1118<=s1118;
Z1119<=s1119;
Z1120<=s1120;
Z1121<=s1121;
Z1122<=s1122;
Z1123<=s1123;
Z1124<=s1124;
Z1125<=s1125;
Z1126<=s1126;
Z1127<=s1127;
Z1128<=s1128;
Z1129<=s1129;
Z1130<=s1130;
Z1131<=s1131;
Z1132<=s1132;
Z1133<=s1133;
Z1134<=s1134;
Z1135<=s1135;
Z1136<=s1136;
Z1137<=s1137;
Z1138<=s1138;
Z1139<=s1139;
Z1140<=s1140;
Z1141<=s1141;
Z1142<=s1142;
Z1143<=s1143;
Z1144<=s1144;
Z1145<=s1145;
Z1146<=s1146;
Z1147<=s1147;
Z1148<=s1148;
Z1149<=s1149;
Z1150<=s1150;
Z1151<=s1151;
Z1152<=s1152;
Z1153<=s1153;
Z1154<=s1154;
Z1155<=s1155;
Z1156<=s1156;
Z1157<=s1157;
Z1158<=s1158;
Z1159<=s1159;
Z1160<=s1160;
Z1161<=s1161;
Z1162<=s1162;
Z1163<=s1163;
Z1164<=s1164;
Z1165<=s1165;
Z1166<=s1166;
Z1167<=s1167;
Z1168<=s1168;
Z1169<=s1169;
Z1170<=s1170;
Z1171<=s1171;
Z1172<=s1172;
Z1173<=s1173;
Z1174<=s1174;
Z1175<=s1175;
Z1176<=s1176;
Z1177<=s1177;
Z1178<=s1178;
Z1179<=s1179;
Z1180<=s1180;
Z1181<=s1181;
Z1182<=s1182;
Z1183<=s1183;
Z1184<=s1184;
Z1185<=s1185;
Z1186<=s1186;
Z1187<=s1187;
Z1188<=s1188;
Z1189<=s1189;
Z1190<=s1190;
Z1191<=s1191;
Z1192<=s1192;
Z1193<=s1193;
Z1194<=s1194;
Z1195<=s1195;
Z1196<=s1196;
Z1197<=s1197;
Z1198<=s1198;
Z1199<=s1199;
Z1200<=s1200;
Z1201<=s1201;
Z1202<=s1202;
Z1203<=s1203;
Z1204<=s1204;
Z1205<=s1205;
Z1206<=s1206;
Z1207<=s1207;
Z1208<=s1208;
Z1209<=s1209;
Z1210<=s1210;
Z1211<=s1211;
Z1212<=s1212;
Z1213<=s1213;
Z1214<=s1214;
Z1215<=s1215;
Z1216<=s1216;
Z1217<=s1217;
Z1218<=s1218;
Z1219<=s1219;
Z1220<=s1220;
Z1221<=s1221;
Z1222<=s1222;
Z1223<=s1223;
Z1224<=s1224;
Z1225<=s1225;
Z1226<=s1226;
Z1227<=s1227;
Z1228<=s1228;
Z1229<=s1229;
Z1230<=s1230;
Z1231<=s1231;
Z1232<=s1232;
Z1233<=s1233;
Z1234<=s1234;
Z1235<=s1235;
Z1236<=s1236;
Z1237<=s1237;
Z1238<=s1238;
Z1239<=s1239;
Z1240<=s1240;
Z1241<=s1241;
Z1242<=s1242;
Z1243<=s1243;
Z1244<=s1244;
Z1245<=s1245;
Z1246<=s1246;
Z1247<=s1247;
Z1248<=s1248;
Z1249<=s1249;
Z1250<=s1250;
Z1251<=s1251;
Z1252<=s1252;
Z1253<=s1253;
Z1254<=s1254;
Z1255<=s1255;
Z1256<=s1256;
Z1257<=s1257;
Z1258<=s1258;
Z1259<=s1259;
Z1260<=s1260;
Z1261<=s1261;
Z1262<=s1262;
Z1263<=s1263;
Z1264<=s1264;
Z1265<=s1265;
Z1266<=s1266;
Z1267<=s1267;
Z1268<=s1268;
Z1269<=s1269;
Z1270<=s1270;
Z1271<=s1271;
Z1272<=s1272;
Z1273<=s1273;
Z1274<=s1274;
Z1275<=s1275;
Z1276<=s1276;
Z1277<=s1277;
Z1278<=s1278;
Z1279<=s1279;
Z1280<=s1280;
Z1281<=s1281;
Z1282<=s1282;
Z1283<=s1283;
Z1284<=s1284;
Z1285<=s1285;
Z1286<=s1286;
Z1287<=s1287;
Z1288<=s1288;
Z1289<=s1289;
Z1290<=s1290;
Z1291<=s1291;
Z1292<=s1292;
Z1293<=s1293;
Z1294<=s1294;
Z1295<=s1295;
Z1296<=s1296;
Z1297<=s1297;
Z1298<=s1298;
Z1299<=s1299;
Z1300<=s1300;
Z1301<=s1301;
Z1302<=s1302;
Z1303<=s1303;
Z1304<=s1304;
Z1305<=s1305;
Z1306<=s1306;
Z1307<=s1307;
Z1308<=s1308;
Z1309<=s1309;
Z1310<=s1310;
Z1311<=s1311;
Z1312<=s1312;
Z1313<=s1313;
Z1314<=s1314;
Z1315<=s1315;
Z1316<=s1316;
Z1317<=s1317;
Z1318<=s1318;
Z1319<=s1319;
Z1320<=s1320;
Z1321<=s1321;
Z1322<=s1322;
Z1323<=s1323;
Z1324<=s1324;
Z1325<=s1325;
Z1326<=s1326;
Z1327<=s1327;
Z1328<=s1328;
Z1329<=s1329;
Z1330<=s1330;
Z1331<=s1331;
Z1332<=s1332;
Z1333<=s1333;
Z1334<=s1334;
Z1335<=s1335;
Z1336<=s1336;
Z1337<=s1337;
Z1338<=s1338;
Z1339<=s1339;
Z1340<=s1340;
Z1341<=s1341;
Z1342<=s1342;
Z1343<=s1343;
Z1344<=s1344;
Z1345<=s1345;
Z1346<=s1346;
Z1347<=s1347;
Z1348<=s1348;
Z1349<=s1349;
Z1350<=s1350;
Z1351<=s1351;
Z1352<=s1352;
Z1353<=s1353;
Z1354<=s1354;
Z1355<=s1355;
Z1356<=s1356;
Z1357<=s1357;
Z1358<=s1358;
Z1359<=s1359;
Z1360<=s1360;
Z1361<=s1361;
Z1362<=s1362;
Z1363<=s1363;
Z1364<=s1364;
Z1365<=s1365;
Z1366<=s1366;
Z1367<=s1367;
Z1368<=s1368;
Z1369<=s1369;
Z1370<=s1370;
Z1371<=s1371;
Z1372<=s1372;
Z1373<=s1373;
Z1374<=s1374;
Z1375<=s1375;
Z1376<=s1376;
Z1377<=s1377;
Z1378<=s1378;
Z1379<=s1379;
Z1380<=s1380;
Z1381<=s1381;
Z1382<=s1382;
Z1383<=s1383;
Z1384<=s1384;
Z1385<=s1385;
Z1386<=s1386;
Z1387<=s1387;
Z1388<=s1388;
Z1389<=s1389;
Z1390<=s1390;
Z1391<=s1391;
Z1392<=s1392;
Z1393<=s1393;
Z1394<=s1394;
Z1395<=s1395;
Z1396<=s1396;
Z1397<=s1397;
Z1398<=s1398;
Z1399<=s1399;
Z1400<=s1400;
Z1401<=s1401;
Z1402<=s1402;
Z1403<=s1403;
Z1404<=s1404;
Z1405<=s1405;
Z1406<=s1406;
Z1407<=s1407;
Z1408<=s1408;
Z1409<=s1409;
Z1410<=s1410;
Z1411<=s1411;
Z1412<=s1412;
Z1413<=s1413;
Z1414<=s1414;
Z1415<=s1415;
Z1416<=s1416;
Z1417<=s1417;
Z1418<=s1418;
Z1419<=s1419;
Z1420<=s1420;
Z1421<=s1421;
Z1422<=s1422;
Z1423<=s1423;
Z1424<=s1424;
Z1425<=s1425;
Z1426<=s1426;
Z1427<=s1427;
Z1428<=s1428;
Z1429<=s1429;
Z1430<=s1430;
Z1431<=s1431;
Z1432<=s1432;
Z1433<=s1433;
Z1434<=s1434;
Z1435<=s1435;
Z1436<=s1436;
Z1437<=s1437;
Z1438<=s1438;
Z1439<=s1439;
Z1440<=s1440;
Z1441<=s1441;
Z1442<=s1442;
Z1443<=s1443;
Z1444<=s1444;
Z1445<=s1445;
Z1446<=s1446;
Z1447<=s1447;
Z1448<=s1448;
Z1449<=s1449;
Z1450<=s1450;
Z1451<=s1451;
Z1452<=s1452;
Z1453<=s1453;
Z1454<=s1454;
Z1455<=s1455;
Z1456<=s1456;
Z1457<=s1457;
Z1458<=s1458;
Z1459<=s1459;
Z1460<=s1460;
Z1461<=s1461;
Z1462<=s1462;
Z1463<=s1463;
Z1464<=s1464;
Z1465<=s1465;
Z1466<=s1466;
Z1467<=s1467;
Z1468<=s1468;
Z1469<=s1469;
Z1470<=s1470;
Z1471<=s1471;
Z1472<=s1472;
Z1473<=s1473;
Z1474<=s1474;
Z1475<=s1475;
Z1476<=s1476;
Z1477<=s1477;
Z1478<=s1478;
Z1479<=s1479;
Z1480<=s1480;
Z1481<=s1481;
Z1482<=s1482;
Z1483<=s1483;
Z1484<=s1484;
Z1485<=s1485;
Z1486<=s1486;
Z1487<=s1487;
Z1488<=s1488;
Z1489<=s1489;
Z1490<=s1490;
Z1491<=s1491;
Z1492<=s1492;
Z1493<=s1493;
Z1494<=s1494;
Z1495<=s1495;
Z1496<=s1496;
Z1497<=s1497;
Z1498<=s1498;
Z1499<=s1499;
Z1500<=s1500;
Z1501<=s1501;
Z1502<=s1502;
Z1503<=s1503;
Z1504<=s1504;
Z1505<=s1505;
Z1506<=s1506;
Z1507<=s1507;
Z1508<=s1508;
Z1509<=s1509;
Z1510<=s1510;
Z1511<=s1511;
Z1512<=s1512;
Z1513<=s1513;
Z1514<=s1514;
Z1515<=s1515;
Z1516<=s1516;
Z1517<=s1517;
Z1518<=s1518;
Z1519<=s1519;
Z1520<=s1520;
Z1521<=s1521;
Z1522<=s1522;
Z1523<=s1523;
Z1524<=s1524;
Z1525<=s1525;
Z1526<=s1526;
Z1527<=s1527;
Z1528<=s1528;
Z1529<=s1529;
Z1530<=s1530;
Z1531<=s1531;
Z1532<=s1532;
Z1533<=s1533;
Z1534<=s1534;
Z1535<=s1535;
Z1536<=s1536;
Z1537<=s1537;
Z1538<=s1538;
Z1539<=s1539;
Z1540<=s1540;
Z1541<=s1541;
Z1542<=s1542;
Z1543<=s1543;
Z1544<=s1544;
Z1545<=s1545;
Z1546<=s1546;
Z1547<=s1547;
Z1548<=s1548;
Z1549<=s1549;
Z1550<=s1550;
Z1551<=s1551;
Z1552<=s1552;
Z1553<=s1553;
Z1554<=s1554;
Z1555<=s1555;
Z1556<=s1556;
Z1557<=s1557;
Z1558<=s1558;
Z1559<=s1559;
Z1560<=s1560;
Z1561<=s1561;
Z1562<=s1562;
Z1563<=s1563;
Z1564<=s1564;
Z1565<=s1565;
Z1566<=s1566;
Z1567<=s1567;
Z1568<=s1568;
Z1569<=s1569;
Z1570<=s1570;
Z1571<=s1571;
Z1572<=s1572;
Z1573<=s1573;
Z1574<=s1574;
Z1575<=s1575;
Z1576<=s1576;
Z1577<=s1577;
Z1578<=s1578;
Z1579<=s1579;
Z1580<=s1580;
Z1581<=s1581;
Z1582<=s1582;
Z1583<=s1583;
Z1584<=s1584;
Z1585<=s1585;
Z1586<=s1586;
Z1587<=s1587;
Z1588<=s1588;
Z1589<=s1589;
Z1590<=s1590;
Z1591<=s1591;
Z1592<=s1592;
Z1593<=s1593;
Z1594<=s1594;
Z1595<=s1595;
Z1596<=s1596;
Z1597<=s1597;
Z1598<=s1598;
Z1599<=s1599;
Z1600<=s1600;
Z1601<=s1601;
Z1602<=s1602;
Z1603<=s1603;
Z1604<=s1604;
Z1605<=s1605;
Z1606<=s1606;
Z1607<=s1607;
Z1608<=s1608;
Z1609<=s1609;
Z1610<=s1610;
Z1611<=s1611;
Z1612<=s1612;
Z1613<=s1613;
Z1614<=s1614;
Z1615<=s1615;
Z1616<=s1616;
Z1617<=s1617;
Z1618<=s1618;
Z1619<=s1619;
Z1620<=s1620;
Z1621<=s1621;
Z1622<=s1622;
Z1623<=s1623;
Z1624<=s1624;
Z1625<=s1625;
Z1626<=s1626;
Z1627<=s1627;
Z1628<=s1628;
Z1629<=s1629;
Z1630<=s1630;
Z1631<=s1631;
Z1632<=s1632;
Z1633<=s1633;
Z1634<=s1634;
Z1635<=s1635;
Z1636<=s1636;
Z1637<=s1637;
Z1638<=s1638;
Z1639<=s1639;
Z1640<=s1640;
Z1641<=s1641;
Z1642<=s1642;
Z1643<=s1643;
Z1644<=s1644;
Z1645<=s1645;
Z1646<=s1646;
Z1647<=s1647;
Z1648<=s1648;
Z1649<=s1649;
Z1650<=s1650;
Z1651<=s1651;
Z1652<=s1652;
Z1653<=s1653;
Z1654<=s1654;
Z1655<=s1655;
Z1656<=s1656;
Z1657<=s1657;
Z1658<=s1658;
Z1659<=s1659;
Z1660<=s1660;
Z1661<=s1661;
Z1662<=s1662;
Z1663<=s1663;
Z1664<=s1664;
Z1665<=s1665;
Z1666<=s1666;
Z1667<=s1667;
Z1668<=s1668;
Z1669<=s1669;
Z1670<=s1670;
Z1671<=s1671;
Z1672<=s1672;
Z1673<=s1673;
Z1674<=s1674;
Z1675<=s1675;
Z1676<=s1676;
Z1677<=s1677;
Z1678<=s1678;
Z1679<=s1679;
Z1680<=s1680;
Z1681<=s1681;
Z1682<=s1682;
Z1683<=s1683;
Z1684<=s1684;
Z1685<=s1685;
Z1686<=s1686;
Z1687<=s1687;
Z1688<=s1688;
Z1689<=s1689;
Z1690<=s1690;
Z1691<=s1691;
Z1692<=s1692;
Z1693<=s1693;
Z1694<=s1694;
Z1695<=s1695;
Z1696<=s1696;
Z1697<=s1697;
Z1698<=s1698;
Z1699<=s1699;
Z1700<=s1700;
Z1701<=s1701;
Z1702<=s1702;
Z1703<=s1703;
Z1704<=s1704;
Z1705<=s1705;
Z1706<=s1706;
Z1707<=s1707;
Z1708<=s1708;
Z1709<=s1709;
Z1710<=s1710;
Z1711<=s1711;
Z1712<=s1712;
Z1713<=s1713;
Z1714<=s1714;
Z1715<=s1715;
Z1716<=s1716;
Z1717<=s1717;
Z1718<=s1718;
Z1719<=s1719;
Z1720<=s1720;
Z1721<=s1721;
Z1722<=s1722;
Z1723<=s1723;
Z1724<=s1724;
Z1725<=s1725;
Z1726<=s1726;
Z1727<=s1727;
Z1728<=s1728;
Z1729<=s1729;
Z1730<=s1730;
Z1731<=s1731;
Z1732<=s1732;
Z1733<=s1733;
Z1734<=s1734;
Z1735<=s1735;
Z1736<=s1736;
Z1737<=s1737;
Z1738<=s1738;
Z1739<=s1739;
Z1740<=s1740;
Z1741<=s1741;
Z1742<=s1742;
Z1743<=s1743;
Z1744<=s1744;
Z1745<=s1745;
Z1746<=s1746;
Z1747<=s1747;
Z1748<=s1748;
Z1749<=s1749;
Z1750<=s1750;
Z1751<=s1751;
Z1752<=s1752;
Z1753<=s1753;
Z1754<=s1754;
Z1755<=s1755;
Z1756<=s1756;
Z1757<=s1757;
Z1758<=s1758;
Z1759<=s1759;
Z1760<=s1760;
Z1761<=s1761;
Z1762<=s1762;
Z1763<=s1763;
Z1764<=s1764;
Z1765<=s1765;
Z1766<=s1766;
Z1767<=s1767;
Z1768<=s1768;
Z1769<=s1769;
Z1770<=s1770;
Z1771<=s1771;
Z1772<=s1772;
Z1773<=s1773;
Z1774<=s1774;
Z1775<=s1775;
Z1776<=s1776;
Z1777<=s1777;
Z1778<=s1778;
Z1779<=s1779;
Z1780<=s1780;
Z1781<=s1781;
Z1782<=s1782;
Z1783<=s1783;
Z1784<=s1784;
Z1785<=s1785;
Z1786<=s1786;
Z1787<=s1787;
Z1788<=s1788;
Z1789<=s1789;
Z1790<=s1790;
Z1791<=s1791;
Z1792<=s1792;
Z1793<=s1793;
Z1794<=s1794;
Z1795<=s1795;
Z1796<=s1796;
Z1797<=s1797;
Z1798<=s1798;
Z1799<=s1799;
Z1800<=s1800;
Z1801<=s1801;
Z1802<=s1802;
Z1803<=s1803;
Z1804<=s1804;
Z1805<=s1805;
Z1806<=s1806;
Z1807<=s1807;
Z1808<=s1808;
Z1809<=s1809;
Z1810<=s1810;
Z1811<=s1811;
Z1812<=s1812;
Z1813<=s1813;
Z1814<=s1814;
Z1815<=s1815;
Z1816<=s1816;
Z1817<=s1817;
Z1818<=s1818;
Z1819<=s1819;
Z1820<=s1820;
Z1821<=s1821;
Z1822<=s1822;
Z1823<=s1823;
Z1824<=s1824;
Z1825<=s1825;
Z1826<=s1826;
Z1827<=s1827;
Z1828<=s1828;
Z1829<=s1829;
Z1830<=s1830;
Z1831<=s1831;
Z1832<=s1832;
Z1833<=s1833;
Z1834<=s1834;
Z1835<=s1835;
Z1836<=s1836;
Z1837<=s1837;
Z1838<=s1838;
Z1839<=s1839;
Z1840<=s1840;
Z1841<=s1841;
Z1842<=s1842;
Z1843<=s1843;
Z1844<=s1844;
Z1845<=s1845;
Z1846<=s1846;
Z1847<=s1847;
Z1848<=s1848;
Z1849<=s1849;
Z1850<=s1850;
Z1851<=s1851;
Z1852<=s1852;
Z1853<=s1853;
Z1854<=s1854;
Z1855<=s1855;
Z1856<=s1856;
Z1857<=s1857;
Z1858<=s1858;
Z1859<=s1859;
Z1860<=s1860;
Z1861<=s1861;
Z1862<=s1862;
Z1863<=s1863;
Z1864<=s1864;
Z1865<=s1865;
Z1866<=s1866;
Z1867<=s1867;
Z1868<=s1868;
Z1869<=s1869;
Z1870<=s1870;
Z1871<=s1871;
Z1872<=s1872;
Z1873<=s1873;
Z1874<=s1874;
Z1875<=s1875;
Z1876<=s1876;
Z1877<=s1877;
Z1878<=s1878;
Z1879<=s1879;
Z1880<=s1880;
Z1881<=s1881;
Z1882<=s1882;
Z1883<=s1883;
Z1884<=s1884;
Z1885<=s1885;
Z1886<=s1886;
Z1887<=s1887;
Z1888<=s1888;
Z1889<=s1889;
Z1890<=s1890;
Z1891<=s1891;
Z1892<=s1892;
Z1893<=s1893;
Z1894<=s1894;
Z1895<=s1895;
Z1896<=s1896;
Z1897<=s1897;
Z1898<=s1898;
Z1899<=s1899;
Z1900<=s1900;
Z1901<=s1901;
Z1902<=s1902;
Z1903<=s1903;
Z1904<=s1904;
Z1905<=s1905;
Z1906<=s1906;
Z1907<=s1907;
Z1908<=s1908;
Z1909<=s1909;
Z1910<=s1910;
Z1911<=s1911;
Z1912<=s1912;
Z1913<=s1913;
Z1914<=s1914;
Z1915<=s1915;
Z1916<=s1916;
Z1917<=s1917;
Z1918<=s1918;
Z1919<=s1919;
Z1920<=s1920;
Z1921<=s1921;
Z1922<=s1922;
Z1923<=s1923;
Z1924<=s1924;
Z1925<=s1925;
Z1926<=s1926;
Z1927<=s1927;
Z1928<=s1928;
Z1929<=s1929;
Z1930<=s1930;
Z1931<=s1931;
Z1932<=s1932;
Z1933<=s1933;
Z1934<=s1934;
Z1935<=s1935;
Z1936<=s1936;
Z1937<=s1937;
Z1938<=s1938;
Z1939<=s1939;
Z1940<=s1940;
Z1941<=s1941;
Z1942<=s1942;
Z1943<=s1943;
Z1944<=s1944;
Z1945<=s1945;
Z1946<=s1946;
Z1947<=s1947;
Z1948<=s1948;
Z1949<=s1949;
Z1950<=s1950;
Z1951<=s1951;
Z1952<=s1952;
Z1953<=s1953;
Z1954<=s1954;
Z1955<=s1955;
Z1956<=s1956;
Z1957<=s1957;
Z1958<=s1958;
Z1959<=s1959;
Z1960<=s1960;
Z1961<=s1961;
Z1962<=s1962;
Z1963<=s1963;
Z1964<=s1964;
Z1965<=s1965;
Z1966<=s1966;
Z1967<=s1967;
Z1968<=s1968;
Z1969<=s1969;
Z1970<=s1970;
Z1971<=s1971;
Z1972<=s1972;
Z1973<=s1973;
Z1974<=s1974;
Z1975<=s1975;
Z1976<=s1976;
Z1977<=s1977;
Z1978<=s1978;
Z1979<=s1979;
Z1980<=s1980;
Z1981<=s1981;
Z1982<=s1982;
Z1983<=s1983;
Z1984<=s1984;
Z1985<=s1985;
Z1986<=s1986;
Z1987<=s1987;
Z1988<=s1988;
Z1989<=s1989;
Z1990<=s1990;
Z1991<=s1991;
Z1992<=s1992;
Z1993<=s1993;
Z1994<=s1994;
Z1995<=s1995;
Z1996<=s1996;
Z1997<=s1997;
Z1998<=s1998;
Z1999<=s1999;
Z2000<=s2000;
Z2001<=s2001;
Z2002<=s2002;
Z2003<=s2003;
Z2004<=s2004;
Z2005<=s2005;
Z2006<=s2006;
Z2007<=s2007;
Z2008<=s2008;
Z2009<=s2009;
Z2010<=s2010;
Z2011<=s2011;
Z2012<=s2012;
Z2013<=s2013;
Z2014<=s2014;
Z2015<=s2015;
Z2016<=s2016;
Z2017<=s2017;
Z2018<=s2018;
Z2019<=s2019;
Z2020<=s2020;
Z2021<=s2021;
Z2022<=s2022;
Z2023<=s2023;
Z2024<=s2024;
Z2025<=s2025;
Z2026<=s2026;
Z2027<=s2027;
Z2028<=s2028;
Z2029<=s2029;
Z2030<=s2030;
Z2031<=s2031;
Z2032<=s2032;
Z2033<=s2033;
Z2034<=s2034;
Z2035<=s2035;
Z2036<=s2036;
Z2037<=s2037;
Z2038<=s2038;
Z2039<=s2039;
Z2040<=s2040;
Z2041<=s2041;
Z2042<=s2042;
Z2043<=s2043;
Z2044<=s2044;
Z2045<=s2045;
Z2046<=s2046;
Z2047<=s2047;
Z2048<=s2048;
Z2049<=s2049;
Z2050<=s2050;
Z2051<=s2051;
Z2052<=s2052;
Z2053<=s2053;
Z2054<=s2054;
Z2055<=s2055;
Z2056<=s2056;
Z2057<=s2057;
Z2058<=s2058;
Z2059<=s2059;
Z2060<=s2060;
Z2061<=s2061;
Z2062<=s2062;
Z2063<=s2063;
Z2064<=s2064;
Z2065<=s2065;
Z2066<=s2066;
Z2067<=s2067;
Z2068<=s2068;
Z2069<=s2069;
Z2070<=s2070;
Z2071<=s2071;
Z2072<=s2072;
Z2073<=s2073;
Z2074<=s2074;
Z2075<=s2075;
Z2076<=s2076;
Z2077<=s2077;
Z2078<=s2078;
Z2079<=s2079;
Z2080<=s2080;
Z2081<=s2081;
Z2082<=s2082;
Z2083<=s2083;
Z2084<=s2084;
Z2085<=s2085;
Z2086<=s2086;
Z2087<=s2087;
Z2088<=s2088;
Z2089<=s2089;
Z2090<=s2090;
Z2091<=s2091;
Z2092<=s2092;
Z2093<=s2093;
Z2094<=s2094;
Z2095<=s2095;
Z2096<=s2096;
Z2097<=s2097;
Z2098<=s2098;
Z2099<=s2099;
Z2100<=s2100;
Z2101<=s2101;
Z2102<=s2102;
Z2103<=s2103;
Z2104<=s2104;
Z2105<=s2105;
Z2106<=s2106;
Z2107<=s2107;
Z2108<=s2108;
Z2109<=s2109;
Z2110<=s2110;
Z2111<=s2111;
Z2112<=s2112;
Z2113<=s2113;
Z2114<=s2114;
Z2115<=s2115;
Z2116<=s2116;
Z2117<=s2117;
Z2118<=s2118;
Z2119<=s2119;
Z2120<=s2120;
Z2121<=s2121;
Z2122<=s2122;
Z2123<=s2123;
Z2124<=s2124;
Z2125<=s2125;
Z2126<=s2126;
Z2127<=s2127;
Z2128<=s2128;
Z2129<=s2129;
Z2130<=s2130;
Z2131<=s2131;
Z2132<=s2132;
Z2133<=s2133;
Z2134<=s2134;
Z2135<=s2135;
Z2136<=s2136;
Z2137<=s2137;
Z2138<=s2138;
Z2139<=s2139;
Z2140<=s2140;
Z2141<=s2141;
Z2142<=s2142;
Z2143<=s2143;
Z2144<=s2144;
Z2145<=s2145;
Z2146<=s2146;
Z2147<=s2147;
Z2148<=s2148;
Z2149<=s2149;
Z2150<=s2150;
Z2151<=s2151;
Z2152<=s2152;
Z2153<=s2153;
Z2154<=s2154;
Z2155<=s2155;
Z2156<=s2156;
Z2157<=s2157;
Z2158<=s2158;
Z2159<=s2159;
Z2160<=s2160;
Z2161<=s2161;
Z2162<=s2162;
Z2163<=s2163;
Z2164<=s2164;
Z2165<=s2165;
Z2166<=s2166;
Z2167<=s2167;
Z2168<=s2168;
Z2169<=s2169;
Z2170<=s2170;
Z2171<=s2171;
Z2172<=s2172;
Z2173<=s2173;
Z2174<=s2174;
Z2175<=s2175;
Z2176<=s2176;
Z2177<=s2177;
Z2178<=s2178;
Z2179<=s2179;
Z2180<=s2180;
Z2181<=s2181;
Z2182<=s2182;
Z2183<=s2183;
Z2184<=s2184;
Z2185<=s2185;
Z2186<=s2186;
Z2187<=s2187;
Z2188<=s2188;
Z2189<=s2189;
Z2190<=s2190;
Z2191<=s2191;
Z2192<=s2192;
Z2193<=s2193;
Z2194<=s2194;
Z2195<=s2195;
Z2196<=s2196;
Z2197<=s2197;
Z2198<=s2198;
Z2199<=s2199;
Z2200<=s2200;
Z2201<=s2201;
Z2202<=s2202;
Z2203<=s2203;
Z2204<=s2204;
Z2205<=s2205;
Z2206<=s2206;
Z2207<=s2207;
Z2208<=s2208;
Z2209<=s2209;
Z2210<=s2210;
Z2211<=s2211;
Z2212<=s2212;
Z2213<=s2213;
Z2214<=s2214;
Z2215<=s2215;
Z2216<=s2216;
Z2217<=s2217;
Z2218<=s2218;
Z2219<=s2219;
Z2220<=s2220;
Z2221<=s2221;
Z2222<=s2222;
Z2223<=s2223;
Z2224<=s2224;
Z2225<=s2225;
Z2226<=s2226;
Z2227<=s2227;
Z2228<=s2228;
Z2229<=s2229;
Z2230<=s2230;
Z2231<=s2231;
Z2232<=s2232;
Z2233<=s2233;
Z2234<=s2234;
Z2235<=s2235;
Z2236<=s2236;
Z2237<=s2237;
Z2238<=s2238;
Z2239<=s2239;
Z2240<=s2240;
Z2241<=s2241;
Z2242<=s2242;
Z2243<=s2243;
Z2244<=s2244;
Z2245<=s2245;
Z2246<=s2246;
Z2247<=s2247;
Z2248<=s2248;
Z2249<=s2249;
Z2250<=s2250;
Z2251<=s2251;
Z2252<=s2252;
Z2253<=s2253;
Z2254<=s2254;
Z2255<=s2255;
Z2256<=s2256;
Z2257<=s2257;
Z2258<=s2258;
Z2259<=s2259;
Z2260<=s2260;
Z2261<=s2261;
Z2262<=s2262;
Z2263<=s2263;
Z2264<=s2264;
Z2265<=s2265;
Z2266<=s2266;
Z2267<=s2267;
Z2268<=s2268;
Z2269<=s2269;
Z2270<=s2270;
Z2271<=s2271;
Z2272<=s2272;
Z2273<=s2273;
Z2274<=s2274;
Z2275<=s2275;
Z2276<=s2276;
Z2277<=s2277;
Z2278<=s2278;
Z2279<=s2279;
Z2280<=s2280;
Z2281<=s2281;
Z2282<=s2282;
Z2283<=s2283;
Z2284<=s2284;
Z2285<=s2285;
Z2286<=s2286;
Z2287<=s2287;
Z2288<=s2288;
Z2289<=s2289;
Z2290<=s2290;
Z2291<=s2291;
Z2292<=s2292;
Z2293<=s2293;
Z2294<=s2294;
Z2295<=s2295;
Z2296<=s2296;
Z2297<=s2297;
Z2298<=s2298;
Z2299<=s2299;
Z2300<=s2300;
Z2301<=s2301;
Z2302<=s2302;
Z2303<=s2303;
Z2304<=s2304;
end;