LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY ldpc IS PORT(
     clk,rst,start_vn,start_cn   :in std_logic;
     Lc1              :in std_logic_vector(8 DOWNTO 0);
     Lc2              :in std_logic_vector(8 DOWNTO 0);
     Lc3              :in std_logic_vector(8 DOWNTO 0);
     Lc4              :in std_logic_vector(8 DOWNTO 0);
     Lc5              :in std_logic_vector(8 DOWNTO 0);
     Lc6              :in std_logic_vector(8 DOWNTO 0);
     Lc7              :in std_logic_vector(8 DOWNTO 0);
     Lc8              :in std_logic_vector(8 DOWNTO 0);
     Lc9              :in std_logic_vector(8 DOWNTO 0);
     Lc10              :in std_logic_vector(8 DOWNTO 0);
     Lc11              :in std_logic_vector(8 DOWNTO 0);
     Lc12              :in std_logic_vector(8 DOWNTO 0);
     Lc13              :in std_logic_vector(8 DOWNTO 0);
     Lc14              :in std_logic_vector(8 DOWNTO 0);
     Lc15              :in std_logic_vector(8 DOWNTO 0);
     Lc16              :in std_logic_vector(8 DOWNTO 0);
     Lc17              :in std_logic_vector(8 DOWNTO 0);
     Lc18              :in std_logic_vector(8 DOWNTO 0);
     Lc19              :in std_logic_vector(8 DOWNTO 0);
     Lc20              :in std_logic_vector(8 DOWNTO 0);
     Lc21              :in std_logic_vector(8 DOWNTO 0);
     Lc22              :in std_logic_vector(8 DOWNTO 0);
     Lc23              :in std_logic_vector(8 DOWNTO 0);
     Lc24              :in std_logic_vector(8 DOWNTO 0);
     Lc25              :in std_logic_vector(8 DOWNTO 0);
     Lc26              :in std_logic_vector(8 DOWNTO 0);
     Lc27              :in std_logic_vector(8 DOWNTO 0);
     Lc28              :in std_logic_vector(8 DOWNTO 0);
     Lc29              :in std_logic_vector(8 DOWNTO 0);
     Lc30              :in std_logic_vector(8 DOWNTO 0);
     Lc31              :in std_logic_vector(8 DOWNTO 0);
     Lc32              :in std_logic_vector(8 DOWNTO 0);
     Lc33              :in std_logic_vector(8 DOWNTO 0);
     Lc34              :in std_logic_vector(8 DOWNTO 0);
     Lc35              :in std_logic_vector(8 DOWNTO 0);
     Lc36              :in std_logic_vector(8 DOWNTO 0);
     Lc37              :in std_logic_vector(8 DOWNTO 0);
     Lc38              :in std_logic_vector(8 DOWNTO 0);
     Lc39              :in std_logic_vector(8 DOWNTO 0);
     Lc40              :in std_logic_vector(8 DOWNTO 0);
     Lc41              :in std_logic_vector(8 DOWNTO 0);
     Lc42              :in std_logic_vector(8 DOWNTO 0);
     Lc43              :in std_logic_vector(8 DOWNTO 0);
     Lc44              :in std_logic_vector(8 DOWNTO 0);
     Lc45              :in std_logic_vector(8 DOWNTO 0);
     Lc46              :in std_logic_vector(8 DOWNTO 0);
     Lc47              :in std_logic_vector(8 DOWNTO 0);
     Lc48              :in std_logic_vector(8 DOWNTO 0);
     Lc49              :in std_logic_vector(8 DOWNTO 0);
     Lc50              :in std_logic_vector(8 DOWNTO 0);
     Lc51              :in std_logic_vector(8 DOWNTO 0);
     Lc52              :in std_logic_vector(8 DOWNTO 0);
     Lc53              :in std_logic_vector(8 DOWNTO 0);
     Lc54              :in std_logic_vector(8 DOWNTO 0);
     Lc55              :in std_logic_vector(8 DOWNTO 0);
     Lc56              :in std_logic_vector(8 DOWNTO 0);
     Lc57              :in std_logic_vector(8 DOWNTO 0);
     Lc58              :in std_logic_vector(8 DOWNTO 0);
     Lc59              :in std_logic_vector(8 DOWNTO 0);
     Lc60              :in std_logic_vector(8 DOWNTO 0);
     Lc61              :in std_logic_vector(8 DOWNTO 0);
     Lc62              :in std_logic_vector(8 DOWNTO 0);
     Lc63              :in std_logic_vector(8 DOWNTO 0);
     Lc64              :in std_logic_vector(8 DOWNTO 0);
     Lc65              :in std_logic_vector(8 DOWNTO 0);
     Lc66              :in std_logic_vector(8 DOWNTO 0);
     Lc67              :in std_logic_vector(8 DOWNTO 0);
     Lc68              :in std_logic_vector(8 DOWNTO 0);
     Lc69              :in std_logic_vector(8 DOWNTO 0);
     Lc70              :in std_logic_vector(8 DOWNTO 0);
     Lc71              :in std_logic_vector(8 DOWNTO 0);
     Lc72              :in std_logic_vector(8 DOWNTO 0);
     Lc73              :in std_logic_vector(8 DOWNTO 0);
     Lc74              :in std_logic_vector(8 DOWNTO 0);
     Lc75              :in std_logic_vector(8 DOWNTO 0);
     Lc76              :in std_logic_vector(8 DOWNTO 0);
     Lc77              :in std_logic_vector(8 DOWNTO 0);
     Lc78              :in std_logic_vector(8 DOWNTO 0);
     Lc79              :in std_logic_vector(8 DOWNTO 0);
     Lc80              :in std_logic_vector(8 DOWNTO 0);
     Lc81              :in std_logic_vector(8 DOWNTO 0);
     Lc82              :in std_logic_vector(8 DOWNTO 0);
     Lc83              :in std_logic_vector(8 DOWNTO 0);
     Lc84              :in std_logic_vector(8 DOWNTO 0);
     Lc85              :in std_logic_vector(8 DOWNTO 0);
     Lc86              :in std_logic_vector(8 DOWNTO 0);
     Lc87              :in std_logic_vector(8 DOWNTO 0);
     Lc88              :in std_logic_vector(8 DOWNTO 0);
     Lc89              :in std_logic_vector(8 DOWNTO 0);
     Lc90              :in std_logic_vector(8 DOWNTO 0);
     Lc91              :in std_logic_vector(8 DOWNTO 0);
     Lc92              :in std_logic_vector(8 DOWNTO 0);
     Lc93              :in std_logic_vector(8 DOWNTO 0);
     Lc94              :in std_logic_vector(8 DOWNTO 0);
     Lc95              :in std_logic_vector(8 DOWNTO 0);
     Lc96              :in std_logic_vector(8 DOWNTO 0);
     Lc97              :in std_logic_vector(8 DOWNTO 0);
     Lc98              :in std_logic_vector(8 DOWNTO 0);
     Lc99              :in std_logic_vector(8 DOWNTO 0);
     Lc100              :in std_logic_vector(8 DOWNTO 0);
     Lc101              :in std_logic_vector(8 DOWNTO 0);
     Lc102              :in std_logic_vector(8 DOWNTO 0);
     Lc103              :in std_logic_vector(8 DOWNTO 0);
     Lc104              :in std_logic_vector(8 DOWNTO 0);
     Lc105              :in std_logic_vector(8 DOWNTO 0);
     Lc106              :in std_logic_vector(8 DOWNTO 0);
     Lc107              :in std_logic_vector(8 DOWNTO 0);
     Lc108              :in std_logic_vector(8 DOWNTO 0);
     Lc109              :in std_logic_vector(8 DOWNTO 0);
     Lc110              :in std_logic_vector(8 DOWNTO 0);
     Lc111              :in std_logic_vector(8 DOWNTO 0);
     Lc112              :in std_logic_vector(8 DOWNTO 0);
     Lc113              :in std_logic_vector(8 DOWNTO 0);
     Lc114              :in std_logic_vector(8 DOWNTO 0);
     Lc115              :in std_logic_vector(8 DOWNTO 0);
     Lc116              :in std_logic_vector(8 DOWNTO 0);
     Lc117              :in std_logic_vector(8 DOWNTO 0);
     Lc118              :in std_logic_vector(8 DOWNTO 0);
     Lc119              :in std_logic_vector(8 DOWNTO 0);
     Lc120              :in std_logic_vector(8 DOWNTO 0);
     Lc121              :in std_logic_vector(8 DOWNTO 0);
     Lc122              :in std_logic_vector(8 DOWNTO 0);
     Lc123              :in std_logic_vector(8 DOWNTO 0);
     Lc124              :in std_logic_vector(8 DOWNTO 0);
     Lc125              :in std_logic_vector(8 DOWNTO 0);
     Lc126              :in std_logic_vector(8 DOWNTO 0);
     Lc127              :in std_logic_vector(8 DOWNTO 0);
     Lc128              :in std_logic_vector(8 DOWNTO 0);
     Lc129              :in std_logic_vector(8 DOWNTO 0);
     Lc130              :in std_logic_vector(8 DOWNTO 0);
     Lc131              :in std_logic_vector(8 DOWNTO 0);
     Lc132              :in std_logic_vector(8 DOWNTO 0);
     Lc133              :in std_logic_vector(8 DOWNTO 0);
     Lc134              :in std_logic_vector(8 DOWNTO 0);
     Lc135              :in std_logic_vector(8 DOWNTO 0);
     Lc136              :in std_logic_vector(8 DOWNTO 0);
     Lc137              :in std_logic_vector(8 DOWNTO 0);
     Lc138              :in std_logic_vector(8 DOWNTO 0);
     Lc139              :in std_logic_vector(8 DOWNTO 0);
     Lc140              :in std_logic_vector(8 DOWNTO 0);
     Lc141              :in std_logic_vector(8 DOWNTO 0);
     Lc142              :in std_logic_vector(8 DOWNTO 0);
     Lc143              :in std_logic_vector(8 DOWNTO 0);
     Lc144              :in std_logic_vector(8 DOWNTO 0);
     Lc145              :in std_logic_vector(8 DOWNTO 0);
     Lc146              :in std_logic_vector(8 DOWNTO 0);
     Lc147              :in std_logic_vector(8 DOWNTO 0);
     Lc148              :in std_logic_vector(8 DOWNTO 0);
     Lc149              :in std_logic_vector(8 DOWNTO 0);
     Lc150              :in std_logic_vector(8 DOWNTO 0);
     Lc151              :in std_logic_vector(8 DOWNTO 0);
     Lc152              :in std_logic_vector(8 DOWNTO 0);
     Lc153              :in std_logic_vector(8 DOWNTO 0);
     Lc154              :in std_logic_vector(8 DOWNTO 0);
     Lc155              :in std_logic_vector(8 DOWNTO 0);
     Lc156              :in std_logic_vector(8 DOWNTO 0);
     Lc157              :in std_logic_vector(8 DOWNTO 0);
     Lc158              :in std_logic_vector(8 DOWNTO 0);
     Lc159              :in std_logic_vector(8 DOWNTO 0);
     Lc160              :in std_logic_vector(8 DOWNTO 0);
     Lc161              :in std_logic_vector(8 DOWNTO 0);
     Lc162              :in std_logic_vector(8 DOWNTO 0);
     Lc163              :in std_logic_vector(8 DOWNTO 0);
     Lc164              :in std_logic_vector(8 DOWNTO 0);
     Lc165              :in std_logic_vector(8 DOWNTO 0);
     Lc166              :in std_logic_vector(8 DOWNTO 0);
     Lc167              :in std_logic_vector(8 DOWNTO 0);
     Lc168              :in std_logic_vector(8 DOWNTO 0);
     Lc169              :in std_logic_vector(8 DOWNTO 0);
     Lc170              :in std_logic_vector(8 DOWNTO 0);
     Lc171              :in std_logic_vector(8 DOWNTO 0);
     Lc172              :in std_logic_vector(8 DOWNTO 0);
     Lc173              :in std_logic_vector(8 DOWNTO 0);
     Lc174              :in std_logic_vector(8 DOWNTO 0);
     Lc175              :in std_logic_vector(8 DOWNTO 0);
     Lc176              :in std_logic_vector(8 DOWNTO 0);
     Lc177              :in std_logic_vector(8 DOWNTO 0);
     Lc178              :in std_logic_vector(8 DOWNTO 0);
     Lc179              :in std_logic_vector(8 DOWNTO 0);
     Lc180              :in std_logic_vector(8 DOWNTO 0);
     Lc181              :in std_logic_vector(8 DOWNTO 0);
     Lc182              :in std_logic_vector(8 DOWNTO 0);
     Lc183              :in std_logic_vector(8 DOWNTO 0);
     Lc184              :in std_logic_vector(8 DOWNTO 0);
     Lc185              :in std_logic_vector(8 DOWNTO 0);
     Lc186              :in std_logic_vector(8 DOWNTO 0);
     Lc187              :in std_logic_vector(8 DOWNTO 0);
     Lc188              :in std_logic_vector(8 DOWNTO 0);
     Lc189              :in std_logic_vector(8 DOWNTO 0);
     Lc190              :in std_logic_vector(8 DOWNTO 0);
     Lc191              :in std_logic_vector(8 DOWNTO 0);
     Lc192              :in std_logic_vector(8 DOWNTO 0);
     Lc193              :in std_logic_vector(8 DOWNTO 0);
     Lc194              :in std_logic_vector(8 DOWNTO 0);
     Lc195              :in std_logic_vector(8 DOWNTO 0);
     Lc196              :in std_logic_vector(8 DOWNTO 0);
     Lc197              :in std_logic_vector(8 DOWNTO 0);
     Lc198              :in std_logic_vector(8 DOWNTO 0);
     Lc199              :in std_logic_vector(8 DOWNTO 0);
     Lc200              :in std_logic_vector(8 DOWNTO 0);
     Lc201              :in std_logic_vector(8 DOWNTO 0);
     Lc202              :in std_logic_vector(8 DOWNTO 0);
     Lc203              :in std_logic_vector(8 DOWNTO 0);
     Lc204              :in std_logic_vector(8 DOWNTO 0);
     Lc205              :in std_logic_vector(8 DOWNTO 0);
     Lc206              :in std_logic_vector(8 DOWNTO 0);
     Lc207              :in std_logic_vector(8 DOWNTO 0);
     Lc208              :in std_logic_vector(8 DOWNTO 0);
     Lc209              :in std_logic_vector(8 DOWNTO 0);
     Lc210              :in std_logic_vector(8 DOWNTO 0);
     Lc211              :in std_logic_vector(8 DOWNTO 0);
     Lc212              :in std_logic_vector(8 DOWNTO 0);
     Lc213              :in std_logic_vector(8 DOWNTO 0);
     Lc214              :in std_logic_vector(8 DOWNTO 0);
     Lc215              :in std_logic_vector(8 DOWNTO 0);
     Lc216              :in std_logic_vector(8 DOWNTO 0);
     Lc217              :in std_logic_vector(8 DOWNTO 0);
     Lc218              :in std_logic_vector(8 DOWNTO 0);
     Lc219              :in std_logic_vector(8 DOWNTO 0);
     Lc220              :in std_logic_vector(8 DOWNTO 0);
     Lc221              :in std_logic_vector(8 DOWNTO 0);
     Lc222              :in std_logic_vector(8 DOWNTO 0);
     Lc223              :in std_logic_vector(8 DOWNTO 0);
     Lc224              :in std_logic_vector(8 DOWNTO 0);
     Lc225              :in std_logic_vector(8 DOWNTO 0);
     Lc226              :in std_logic_vector(8 DOWNTO 0);
     Lc227              :in std_logic_vector(8 DOWNTO 0);
     Lc228              :in std_logic_vector(8 DOWNTO 0);
     Lc229              :in std_logic_vector(8 DOWNTO 0);
     Lc230              :in std_logic_vector(8 DOWNTO 0);
     Lc231              :in std_logic_vector(8 DOWNTO 0);
     Lc232              :in std_logic_vector(8 DOWNTO 0);
     Lc233              :in std_logic_vector(8 DOWNTO 0);
     Lc234              :in std_logic_vector(8 DOWNTO 0);
     Lc235              :in std_logic_vector(8 DOWNTO 0);
     Lc236              :in std_logic_vector(8 DOWNTO 0);
     Lc237              :in std_logic_vector(8 DOWNTO 0);
     Lc238              :in std_logic_vector(8 DOWNTO 0);
     Lc239              :in std_logic_vector(8 DOWNTO 0);
     Lc240              :in std_logic_vector(8 DOWNTO 0);
     Lc241              :in std_logic_vector(8 DOWNTO 0);
     Lc242              :in std_logic_vector(8 DOWNTO 0);
     Lc243              :in std_logic_vector(8 DOWNTO 0);
     Lc244              :in std_logic_vector(8 DOWNTO 0);
     Lc245              :in std_logic_vector(8 DOWNTO 0);
     Lc246              :in std_logic_vector(8 DOWNTO 0);
     Lc247              :in std_logic_vector(8 DOWNTO 0);
     Lc248              :in std_logic_vector(8 DOWNTO 0);
     Lc249              :in std_logic_vector(8 DOWNTO 0);
     Lc250              :in std_logic_vector(8 DOWNTO 0);
     Lc251              :in std_logic_vector(8 DOWNTO 0);
     Lc252              :in std_logic_vector(8 DOWNTO 0);
     Lc253              :in std_logic_vector(8 DOWNTO 0);
     Lc254              :in std_logic_vector(8 DOWNTO 0);
     Lc255              :in std_logic_vector(8 DOWNTO 0);
     Lc256              :in std_logic_vector(8 DOWNTO 0);
     Lc257              :in std_logic_vector(8 DOWNTO 0);
     Lc258              :in std_logic_vector(8 DOWNTO 0);
     Lc259              :in std_logic_vector(8 DOWNTO 0);
     Lc260              :in std_logic_vector(8 DOWNTO 0);
     Lc261              :in std_logic_vector(8 DOWNTO 0);
     Lc262              :in std_logic_vector(8 DOWNTO 0);
     Lc263              :in std_logic_vector(8 DOWNTO 0);
     Lc264              :in std_logic_vector(8 DOWNTO 0);
     Lc265              :in std_logic_vector(8 DOWNTO 0);
     Lc266              :in std_logic_vector(8 DOWNTO 0);
     Lc267              :in std_logic_vector(8 DOWNTO 0);
     Lc268              :in std_logic_vector(8 DOWNTO 0);
     Lc269              :in std_logic_vector(8 DOWNTO 0);
     Lc270              :in std_logic_vector(8 DOWNTO 0);
     Lc271              :in std_logic_vector(8 DOWNTO 0);
     Lc272              :in std_logic_vector(8 DOWNTO 0);
     Lc273              :in std_logic_vector(8 DOWNTO 0);
     Lc274              :in std_logic_vector(8 DOWNTO 0);
     Lc275              :in std_logic_vector(8 DOWNTO 0);
     Lc276              :in std_logic_vector(8 DOWNTO 0);
     Lc277              :in std_logic_vector(8 DOWNTO 0);
     Lc278              :in std_logic_vector(8 DOWNTO 0);
     Lc279              :in std_logic_vector(8 DOWNTO 0);
     Lc280              :in std_logic_vector(8 DOWNTO 0);
     Lc281              :in std_logic_vector(8 DOWNTO 0);
     Lc282              :in std_logic_vector(8 DOWNTO 0);
     Lc283              :in std_logic_vector(8 DOWNTO 0);
     Lc284              :in std_logic_vector(8 DOWNTO 0);
     Lc285              :in std_logic_vector(8 DOWNTO 0);
     Lc286              :in std_logic_vector(8 DOWNTO 0);
     Lc287              :in std_logic_vector(8 DOWNTO 0);
     Lc288              :in std_logic_vector(8 DOWNTO 0);
     Lc289              :in std_logic_vector(8 DOWNTO 0);
     Lc290              :in std_logic_vector(8 DOWNTO 0);
     Lc291              :in std_logic_vector(8 DOWNTO 0);
     Lc292              :in std_logic_vector(8 DOWNTO 0);
     Lc293              :in std_logic_vector(8 DOWNTO 0);
     Lc294              :in std_logic_vector(8 DOWNTO 0);
     Lc295              :in std_logic_vector(8 DOWNTO 0);
     Lc296              :in std_logic_vector(8 DOWNTO 0);
     Lc297              :in std_logic_vector(8 DOWNTO 0);
     Lc298              :in std_logic_vector(8 DOWNTO 0);
     Lc299              :in std_logic_vector(8 DOWNTO 0);
     Lc300              :in std_logic_vector(8 DOWNTO 0);
     Lc301              :in std_logic_vector(8 DOWNTO 0);
     Lc302              :in std_logic_vector(8 DOWNTO 0);
     Lc303              :in std_logic_vector(8 DOWNTO 0);
     Lc304              :in std_logic_vector(8 DOWNTO 0);
     Lc305              :in std_logic_vector(8 DOWNTO 0);
     Lc306              :in std_logic_vector(8 DOWNTO 0);
     Lc307              :in std_logic_vector(8 DOWNTO 0);
     Lc308              :in std_logic_vector(8 DOWNTO 0);
     Lc309              :in std_logic_vector(8 DOWNTO 0);
     Lc310              :in std_logic_vector(8 DOWNTO 0);
     Lc311              :in std_logic_vector(8 DOWNTO 0);
     Lc312              :in std_logic_vector(8 DOWNTO 0);
     Lc313              :in std_logic_vector(8 DOWNTO 0);
     Lc314              :in std_logic_vector(8 DOWNTO 0);
     Lc315              :in std_logic_vector(8 DOWNTO 0);
     Lc316              :in std_logic_vector(8 DOWNTO 0);
     Lc317              :in std_logic_vector(8 DOWNTO 0);
     Lc318              :in std_logic_vector(8 DOWNTO 0);
     Lc319              :in std_logic_vector(8 DOWNTO 0);
     Lc320              :in std_logic_vector(8 DOWNTO 0);
     Lc321              :in std_logic_vector(8 DOWNTO 0);
     Lc322              :in std_logic_vector(8 DOWNTO 0);
     Lc323              :in std_logic_vector(8 DOWNTO 0);
     Lc324              :in std_logic_vector(8 DOWNTO 0);
     Lc325              :in std_logic_vector(8 DOWNTO 0);
     Lc326              :in std_logic_vector(8 DOWNTO 0);
     Lc327              :in std_logic_vector(8 DOWNTO 0);
     Lc328              :in std_logic_vector(8 DOWNTO 0);
     Lc329              :in std_logic_vector(8 DOWNTO 0);
     Lc330              :in std_logic_vector(8 DOWNTO 0);
     Lc331              :in std_logic_vector(8 DOWNTO 0);
     Lc332              :in std_logic_vector(8 DOWNTO 0);
     Lc333              :in std_logic_vector(8 DOWNTO 0);
     Lc334              :in std_logic_vector(8 DOWNTO 0);
     Lc335              :in std_logic_vector(8 DOWNTO 0);
     Lc336              :in std_logic_vector(8 DOWNTO 0);
     Lc337              :in std_logic_vector(8 DOWNTO 0);
     Lc338              :in std_logic_vector(8 DOWNTO 0);
     Lc339              :in std_logic_vector(8 DOWNTO 0);
     Lc340              :in std_logic_vector(8 DOWNTO 0);
     Lc341              :in std_logic_vector(8 DOWNTO 0);
     Lc342              :in std_logic_vector(8 DOWNTO 0);
     Lc343              :in std_logic_vector(8 DOWNTO 0);
     Lc344              :in std_logic_vector(8 DOWNTO 0);
     Lc345              :in std_logic_vector(8 DOWNTO 0);
     Lc346              :in std_logic_vector(8 DOWNTO 0);
     Lc347              :in std_logic_vector(8 DOWNTO 0);
     Lc348              :in std_logic_vector(8 DOWNTO 0);
     Lc349              :in std_logic_vector(8 DOWNTO 0);
     Lc350              :in std_logic_vector(8 DOWNTO 0);
     Lc351              :in std_logic_vector(8 DOWNTO 0);
     Lc352              :in std_logic_vector(8 DOWNTO 0);
     Lc353              :in std_logic_vector(8 DOWNTO 0);
     Lc354              :in std_logic_vector(8 DOWNTO 0);
     Lc355              :in std_logic_vector(8 DOWNTO 0);
     Lc356              :in std_logic_vector(8 DOWNTO 0);
     Lc357              :in std_logic_vector(8 DOWNTO 0);
     Lc358              :in std_logic_vector(8 DOWNTO 0);
     Lc359              :in std_logic_vector(8 DOWNTO 0);
     Lc360              :in std_logic_vector(8 DOWNTO 0);
     Lc361              :in std_logic_vector(8 DOWNTO 0);
     Lc362              :in std_logic_vector(8 DOWNTO 0);
     Lc363              :in std_logic_vector(8 DOWNTO 0);
     Lc364              :in std_logic_vector(8 DOWNTO 0);
     Lc365              :in std_logic_vector(8 DOWNTO 0);
     Lc366              :in std_logic_vector(8 DOWNTO 0);
     Lc367              :in std_logic_vector(8 DOWNTO 0);
     Lc368              :in std_logic_vector(8 DOWNTO 0);
     Lc369              :in std_logic_vector(8 DOWNTO 0);
     Lc370              :in std_logic_vector(8 DOWNTO 0);
     Lc371              :in std_logic_vector(8 DOWNTO 0);
     Lc372              :in std_logic_vector(8 DOWNTO 0);
     Lc373              :in std_logic_vector(8 DOWNTO 0);
     Lc374              :in std_logic_vector(8 DOWNTO 0);
     Lc375              :in std_logic_vector(8 DOWNTO 0);
     Lc376              :in std_logic_vector(8 DOWNTO 0);
     Lc377              :in std_logic_vector(8 DOWNTO 0);
     Lc378              :in std_logic_vector(8 DOWNTO 0);
     Lc379              :in std_logic_vector(8 DOWNTO 0);
     Lc380              :in std_logic_vector(8 DOWNTO 0);
     Lc381              :in std_logic_vector(8 DOWNTO 0);
     Lc382              :in std_logic_vector(8 DOWNTO 0);
     Lc383              :in std_logic_vector(8 DOWNTO 0);
     Lc384              :in std_logic_vector(8 DOWNTO 0);
     Lc385              :in std_logic_vector(8 DOWNTO 0);
     Lc386              :in std_logic_vector(8 DOWNTO 0);
     Lc387              :in std_logic_vector(8 DOWNTO 0);
     Lc388              :in std_logic_vector(8 DOWNTO 0);
     Lc389              :in std_logic_vector(8 DOWNTO 0);
     Lc390              :in std_logic_vector(8 DOWNTO 0);
     Lc391              :in std_logic_vector(8 DOWNTO 0);
     Lc392              :in std_logic_vector(8 DOWNTO 0);
     Lc393              :in std_logic_vector(8 DOWNTO 0);
     Lc394              :in std_logic_vector(8 DOWNTO 0);
     Lc395              :in std_logic_vector(8 DOWNTO 0);
     Lc396              :in std_logic_vector(8 DOWNTO 0);
     Lc397              :in std_logic_vector(8 DOWNTO 0);
     Lc398              :in std_logic_vector(8 DOWNTO 0);
     Lc399              :in std_logic_vector(8 DOWNTO 0);
     Lc400              :in std_logic_vector(8 DOWNTO 0);
     Lc401              :in std_logic_vector(8 DOWNTO 0);
     Lc402              :in std_logic_vector(8 DOWNTO 0);
     Lc403              :in std_logic_vector(8 DOWNTO 0);
     Lc404              :in std_logic_vector(8 DOWNTO 0);
     Lc405              :in std_logic_vector(8 DOWNTO 0);
     Lc406              :in std_logic_vector(8 DOWNTO 0);
     Lc407              :in std_logic_vector(8 DOWNTO 0);
     Lc408              :in std_logic_vector(8 DOWNTO 0);
     Lc409              :in std_logic_vector(8 DOWNTO 0);
     Lc410              :in std_logic_vector(8 DOWNTO 0);
     Lc411              :in std_logic_vector(8 DOWNTO 0);
     Lc412              :in std_logic_vector(8 DOWNTO 0);
     Lc413              :in std_logic_vector(8 DOWNTO 0);
     Lc414              :in std_logic_vector(8 DOWNTO 0);
     Lc415              :in std_logic_vector(8 DOWNTO 0);
     Lc416              :in std_logic_vector(8 DOWNTO 0);
     Lc417              :in std_logic_vector(8 DOWNTO 0);
     Lc418              :in std_logic_vector(8 DOWNTO 0);
     Lc419              :in std_logic_vector(8 DOWNTO 0);
     Lc420              :in std_logic_vector(8 DOWNTO 0);
     Lc421              :in std_logic_vector(8 DOWNTO 0);
     Lc422              :in std_logic_vector(8 DOWNTO 0);
     Lc423              :in std_logic_vector(8 DOWNTO 0);
     Lc424              :in std_logic_vector(8 DOWNTO 0);
     Lc425              :in std_logic_vector(8 DOWNTO 0);
     Lc426              :in std_logic_vector(8 DOWNTO 0);
     Lc427              :in std_logic_vector(8 DOWNTO 0);
     Lc428              :in std_logic_vector(8 DOWNTO 0);
     Lc429              :in std_logic_vector(8 DOWNTO 0);
     Lc430              :in std_logic_vector(8 DOWNTO 0);
     Lc431              :in std_logic_vector(8 DOWNTO 0);
     Lc432              :in std_logic_vector(8 DOWNTO 0);
     Lc433              :in std_logic_vector(8 DOWNTO 0);
     Lc434              :in std_logic_vector(8 DOWNTO 0);
     Lc435              :in std_logic_vector(8 DOWNTO 0);
     Lc436              :in std_logic_vector(8 DOWNTO 0);
     Lc437              :in std_logic_vector(8 DOWNTO 0);
     Lc438              :in std_logic_vector(8 DOWNTO 0);
     Lc439              :in std_logic_vector(8 DOWNTO 0);
     Lc440              :in std_logic_vector(8 DOWNTO 0);
     Lc441              :in std_logic_vector(8 DOWNTO 0);
     Lc442              :in std_logic_vector(8 DOWNTO 0);
     Lc443              :in std_logic_vector(8 DOWNTO 0);
     Lc444              :in std_logic_vector(8 DOWNTO 0);
     Lc445              :in std_logic_vector(8 DOWNTO 0);
     Lc446              :in std_logic_vector(8 DOWNTO 0);
     Lc447              :in std_logic_vector(8 DOWNTO 0);
     Lc448              :in std_logic_vector(8 DOWNTO 0);
     Lc449              :in std_logic_vector(8 DOWNTO 0);
     Lc450              :in std_logic_vector(8 DOWNTO 0);
     Lc451              :in std_logic_vector(8 DOWNTO 0);
     Lc452              :in std_logic_vector(8 DOWNTO 0);
     Lc453              :in std_logic_vector(8 DOWNTO 0);
     Lc454              :in std_logic_vector(8 DOWNTO 0);
     Lc455              :in std_logic_vector(8 DOWNTO 0);
     Lc456              :in std_logic_vector(8 DOWNTO 0);
     Lc457              :in std_logic_vector(8 DOWNTO 0);
     Lc458              :in std_logic_vector(8 DOWNTO 0);
     Lc459              :in std_logic_vector(8 DOWNTO 0);
     Lc460              :in std_logic_vector(8 DOWNTO 0);
     Lc461              :in std_logic_vector(8 DOWNTO 0);
     Lc462              :in std_logic_vector(8 DOWNTO 0);
     Lc463              :in std_logic_vector(8 DOWNTO 0);
     Lc464              :in std_logic_vector(8 DOWNTO 0);
     Lc465              :in std_logic_vector(8 DOWNTO 0);
     Lc466              :in std_logic_vector(8 DOWNTO 0);
     Lc467              :in std_logic_vector(8 DOWNTO 0);
     Lc468              :in std_logic_vector(8 DOWNTO 0);
     Lc469              :in std_logic_vector(8 DOWNTO 0);
     Lc470              :in std_logic_vector(8 DOWNTO 0);
     Lc471              :in std_logic_vector(8 DOWNTO 0);
     Lc472              :in std_logic_vector(8 DOWNTO 0);
     Lc473              :in std_logic_vector(8 DOWNTO 0);
     Lc474              :in std_logic_vector(8 DOWNTO 0);
     Lc475              :in std_logic_vector(8 DOWNTO 0);
     Lc476              :in std_logic_vector(8 DOWNTO 0);
     Lc477              :in std_logic_vector(8 DOWNTO 0);
     Lc478              :in std_logic_vector(8 DOWNTO 0);
     Lc479              :in std_logic_vector(8 DOWNTO 0);
     Lc480              :in std_logic_vector(8 DOWNTO 0);
     Lc481              :in std_logic_vector(8 DOWNTO 0);
     Lc482              :in std_logic_vector(8 DOWNTO 0);
     Lc483              :in std_logic_vector(8 DOWNTO 0);
     Lc484              :in std_logic_vector(8 DOWNTO 0);
     Lc485              :in std_logic_vector(8 DOWNTO 0);
     Lc486              :in std_logic_vector(8 DOWNTO 0);
     Lc487              :in std_logic_vector(8 DOWNTO 0);
     Lc488              :in std_logic_vector(8 DOWNTO 0);
     Lc489              :in std_logic_vector(8 DOWNTO 0);
     Lc490              :in std_logic_vector(8 DOWNTO 0);
     Lc491              :in std_logic_vector(8 DOWNTO 0);
     Lc492              :in std_logic_vector(8 DOWNTO 0);
     Lc493              :in std_logic_vector(8 DOWNTO 0);
     Lc494              :in std_logic_vector(8 DOWNTO 0);
     Lc495              :in std_logic_vector(8 DOWNTO 0);
     Lc496              :in std_logic_vector(8 DOWNTO 0);
     Lc497              :in std_logic_vector(8 DOWNTO 0);
     Lc498              :in std_logic_vector(8 DOWNTO 0);
     Lc499              :in std_logic_vector(8 DOWNTO 0);
     Lc500              :in std_logic_vector(8 DOWNTO 0);
     Lc501              :in std_logic_vector(8 DOWNTO 0);
     Lc502              :in std_logic_vector(8 DOWNTO 0);
     Lc503              :in std_logic_vector(8 DOWNTO 0);
     Lc504              :in std_logic_vector(8 DOWNTO 0);
     Lc505              :in std_logic_vector(8 DOWNTO 0);
     Lc506              :in std_logic_vector(8 DOWNTO 0);
     Lc507              :in std_logic_vector(8 DOWNTO 0);
     Lc508              :in std_logic_vector(8 DOWNTO 0);
     Lc509              :in std_logic_vector(8 DOWNTO 0);
     Lc510              :in std_logic_vector(8 DOWNTO 0);
     Lc511              :in std_logic_vector(8 DOWNTO 0);
     Lc512              :in std_logic_vector(8 DOWNTO 0);
     Lc513              :in std_logic_vector(8 DOWNTO 0);
     Lc514              :in std_logic_vector(8 DOWNTO 0);
     Lc515              :in std_logic_vector(8 DOWNTO 0);
     Lc516              :in std_logic_vector(8 DOWNTO 0);
     Lc517              :in std_logic_vector(8 DOWNTO 0);
     Lc518              :in std_logic_vector(8 DOWNTO 0);
     Lc519              :in std_logic_vector(8 DOWNTO 0);
     Lc520              :in std_logic_vector(8 DOWNTO 0);
     Lc521              :in std_logic_vector(8 DOWNTO 0);
     Lc522              :in std_logic_vector(8 DOWNTO 0);
     Lc523              :in std_logic_vector(8 DOWNTO 0);
     Lc524              :in std_logic_vector(8 DOWNTO 0);
     Lc525              :in std_logic_vector(8 DOWNTO 0);
     Lc526              :in std_logic_vector(8 DOWNTO 0);
     Lc527              :in std_logic_vector(8 DOWNTO 0);
     Lc528              :in std_logic_vector(8 DOWNTO 0);
     Lc529              :in std_logic_vector(8 DOWNTO 0);
     Lc530              :in std_logic_vector(8 DOWNTO 0);
     Lc531              :in std_logic_vector(8 DOWNTO 0);
     Lc532              :in std_logic_vector(8 DOWNTO 0);
     Lc533              :in std_logic_vector(8 DOWNTO 0);
     Lc534              :in std_logic_vector(8 DOWNTO 0);
     Lc535              :in std_logic_vector(8 DOWNTO 0);
     Lc536              :in std_logic_vector(8 DOWNTO 0);
     Lc537              :in std_logic_vector(8 DOWNTO 0);
     Lc538              :in std_logic_vector(8 DOWNTO 0);
     Lc539              :in std_logic_vector(8 DOWNTO 0);
     Lc540              :in std_logic_vector(8 DOWNTO 0);
     Lc541              :in std_logic_vector(8 DOWNTO 0);
     Lc542              :in std_logic_vector(8 DOWNTO 0);
     Lc543              :in std_logic_vector(8 DOWNTO 0);
     Lc544              :in std_logic_vector(8 DOWNTO 0);
     Lc545              :in std_logic_vector(8 DOWNTO 0);
     Lc546              :in std_logic_vector(8 DOWNTO 0);
     Lc547              :in std_logic_vector(8 DOWNTO 0);
     Lc548              :in std_logic_vector(8 DOWNTO 0);
     Lc549              :in std_logic_vector(8 DOWNTO 0);
     Lc550              :in std_logic_vector(8 DOWNTO 0);
     Lc551              :in std_logic_vector(8 DOWNTO 0);
     Lc552              :in std_logic_vector(8 DOWNTO 0);
     Lc553              :in std_logic_vector(8 DOWNTO 0);
     Lc554              :in std_logic_vector(8 DOWNTO 0);
     Lc555              :in std_logic_vector(8 DOWNTO 0);
     Lc556              :in std_logic_vector(8 DOWNTO 0);
     Lc557              :in std_logic_vector(8 DOWNTO 0);
     Lc558              :in std_logic_vector(8 DOWNTO 0);
     Lc559              :in std_logic_vector(8 DOWNTO 0);
     Lc560              :in std_logic_vector(8 DOWNTO 0);
     Lc561              :in std_logic_vector(8 DOWNTO 0);
     Lc562              :in std_logic_vector(8 DOWNTO 0);
     Lc563              :in std_logic_vector(8 DOWNTO 0);
     Lc564              :in std_logic_vector(8 DOWNTO 0);
     Lc565              :in std_logic_vector(8 DOWNTO 0);
     Lc566              :in std_logic_vector(8 DOWNTO 0);
     Lc567              :in std_logic_vector(8 DOWNTO 0);
     Lc568              :in std_logic_vector(8 DOWNTO 0);
     Lc569              :in std_logic_vector(8 DOWNTO 0);
     Lc570              :in std_logic_vector(8 DOWNTO 0);
     Lc571              :in std_logic_vector(8 DOWNTO 0);
     Lc572              :in std_logic_vector(8 DOWNTO 0);
     Lc573              :in std_logic_vector(8 DOWNTO 0);
     Lc574              :in std_logic_vector(8 DOWNTO 0);
     Lc575              :in std_logic_vector(8 DOWNTO 0);
     Lc576              :in std_logic_vector(8 DOWNTO 0);
     Lc577              :in std_logic_vector(8 DOWNTO 0);
     Lc578              :in std_logic_vector(8 DOWNTO 0);
     Lc579              :in std_logic_vector(8 DOWNTO 0);
     Lc580              :in std_logic_vector(8 DOWNTO 0);
     Lc581              :in std_logic_vector(8 DOWNTO 0);
     Lc582              :in std_logic_vector(8 DOWNTO 0);
     Lc583              :in std_logic_vector(8 DOWNTO 0);
     Lc584              :in std_logic_vector(8 DOWNTO 0);
     Lc585              :in std_logic_vector(8 DOWNTO 0);
     Lc586              :in std_logic_vector(8 DOWNTO 0);
     Lc587              :in std_logic_vector(8 DOWNTO 0);
     Lc588              :in std_logic_vector(8 DOWNTO 0);
     Lc589              :in std_logic_vector(8 DOWNTO 0);
     Lc590              :in std_logic_vector(8 DOWNTO 0);
     Lc591              :in std_logic_vector(8 DOWNTO 0);
     Lc592              :in std_logic_vector(8 DOWNTO 0);
     Lc593              :in std_logic_vector(8 DOWNTO 0);
     Lc594              :in std_logic_vector(8 DOWNTO 0);
     Lc595              :in std_logic_vector(8 DOWNTO 0);
     Lc596              :in std_logic_vector(8 DOWNTO 0);
     Lc597              :in std_logic_vector(8 DOWNTO 0);
     Lc598              :in std_logic_vector(8 DOWNTO 0);
     Lc599              :in std_logic_vector(8 DOWNTO 0);
     Lc600              :in std_logic_vector(8 DOWNTO 0);
     Lc601              :in std_logic_vector(8 DOWNTO 0);
     Lc602              :in std_logic_vector(8 DOWNTO 0);
     Lc603              :in std_logic_vector(8 DOWNTO 0);
     Lc604              :in std_logic_vector(8 DOWNTO 0);
     Lc605              :in std_logic_vector(8 DOWNTO 0);
     Lc606              :in std_logic_vector(8 DOWNTO 0);
     Lc607              :in std_logic_vector(8 DOWNTO 0);
     Lc608              :in std_logic_vector(8 DOWNTO 0);
     Lc609              :in std_logic_vector(8 DOWNTO 0);
     Lc610              :in std_logic_vector(8 DOWNTO 0);
     Lc611              :in std_logic_vector(8 DOWNTO 0);
     Lc612              :in std_logic_vector(8 DOWNTO 0);
     Lc613              :in std_logic_vector(8 DOWNTO 0);
     Lc614              :in std_logic_vector(8 DOWNTO 0);
     Lc615              :in std_logic_vector(8 DOWNTO 0);
     Lc616              :in std_logic_vector(8 DOWNTO 0);
     Lc617              :in std_logic_vector(8 DOWNTO 0);
     Lc618              :in std_logic_vector(8 DOWNTO 0);
     Lc619              :in std_logic_vector(8 DOWNTO 0);
     Lc620              :in std_logic_vector(8 DOWNTO 0);
     Lc621              :in std_logic_vector(8 DOWNTO 0);
     Lc622              :in std_logic_vector(8 DOWNTO 0);
     Lc623              :in std_logic_vector(8 DOWNTO 0);
     Lc624              :in std_logic_vector(8 DOWNTO 0);
     Lc625              :in std_logic_vector(8 DOWNTO 0);
     Lc626              :in std_logic_vector(8 DOWNTO 0);
     Lc627              :in std_logic_vector(8 DOWNTO 0);
     Lc628              :in std_logic_vector(8 DOWNTO 0);
     Lc629              :in std_logic_vector(8 DOWNTO 0);
     Lc630              :in std_logic_vector(8 DOWNTO 0);
     Lc631              :in std_logic_vector(8 DOWNTO 0);
     Lc632              :in std_logic_vector(8 DOWNTO 0);
     Lc633              :in std_logic_vector(8 DOWNTO 0);
     Lc634              :in std_logic_vector(8 DOWNTO 0);
     Lc635              :in std_logic_vector(8 DOWNTO 0);
     Lc636              :in std_logic_vector(8 DOWNTO 0);
     Lc637              :in std_logic_vector(8 DOWNTO 0);
     Lc638              :in std_logic_vector(8 DOWNTO 0);
     Lc639              :in std_logic_vector(8 DOWNTO 0);
     Lc640              :in std_logic_vector(8 DOWNTO 0);
     Lc641              :in std_logic_vector(8 DOWNTO 0);
     Lc642              :in std_logic_vector(8 DOWNTO 0);
     Lc643              :in std_logic_vector(8 DOWNTO 0);
     Lc644              :in std_logic_vector(8 DOWNTO 0);
     Lc645              :in std_logic_vector(8 DOWNTO 0);
     Lc646              :in std_logic_vector(8 DOWNTO 0);
     Lc647              :in std_logic_vector(8 DOWNTO 0);
     Lc648              :in std_logic_vector(8 DOWNTO 0);
     Lc649              :in std_logic_vector(8 DOWNTO 0);
     Lc650              :in std_logic_vector(8 DOWNTO 0);
     Lc651              :in std_logic_vector(8 DOWNTO 0);
     Lc652              :in std_logic_vector(8 DOWNTO 0);
     Lc653              :in std_logic_vector(8 DOWNTO 0);
     Lc654              :in std_logic_vector(8 DOWNTO 0);
     Lc655              :in std_logic_vector(8 DOWNTO 0);
     Lc656              :in std_logic_vector(8 DOWNTO 0);
     Lc657              :in std_logic_vector(8 DOWNTO 0);
     Lc658              :in std_logic_vector(8 DOWNTO 0);
     Lc659              :in std_logic_vector(8 DOWNTO 0);
     Lc660              :in std_logic_vector(8 DOWNTO 0);
     Lc661              :in std_logic_vector(8 DOWNTO 0);
     Lc662              :in std_logic_vector(8 DOWNTO 0);
     Lc663              :in std_logic_vector(8 DOWNTO 0);
     Lc664              :in std_logic_vector(8 DOWNTO 0);
     Lc665              :in std_logic_vector(8 DOWNTO 0);
     Lc666              :in std_logic_vector(8 DOWNTO 0);
     Lc667              :in std_logic_vector(8 DOWNTO 0);
     Lc668              :in std_logic_vector(8 DOWNTO 0);
     Lc669              :in std_logic_vector(8 DOWNTO 0);
     Lc670              :in std_logic_vector(8 DOWNTO 0);
     Lc671              :in std_logic_vector(8 DOWNTO 0);
     Lc672              :in std_logic_vector(8 DOWNTO 0);
     Lc673              :in std_logic_vector(8 DOWNTO 0);
     Lc674              :in std_logic_vector(8 DOWNTO 0);
     Lc675              :in std_logic_vector(8 DOWNTO 0);
     Lc676              :in std_logic_vector(8 DOWNTO 0);
     Lc677              :in std_logic_vector(8 DOWNTO 0);
     Lc678              :in std_logic_vector(8 DOWNTO 0);
     Lc679              :in std_logic_vector(8 DOWNTO 0);
     Lc680              :in std_logic_vector(8 DOWNTO 0);
     Lc681              :in std_logic_vector(8 DOWNTO 0);
     Lc682              :in std_logic_vector(8 DOWNTO 0);
     Lc683              :in std_logic_vector(8 DOWNTO 0);
     Lc684              :in std_logic_vector(8 DOWNTO 0);
     Lc685              :in std_logic_vector(8 DOWNTO 0);
     Lc686              :in std_logic_vector(8 DOWNTO 0);
     Lc687              :in std_logic_vector(8 DOWNTO 0);
     Lc688              :in std_logic_vector(8 DOWNTO 0);
     Lc689              :in std_logic_vector(8 DOWNTO 0);
     Lc690              :in std_logic_vector(8 DOWNTO 0);
     Lc691              :in std_logic_vector(8 DOWNTO 0);
     Lc692              :in std_logic_vector(8 DOWNTO 0);
     Lc693              :in std_logic_vector(8 DOWNTO 0);
     Lc694              :in std_logic_vector(8 DOWNTO 0);
     Lc695              :in std_logic_vector(8 DOWNTO 0);
     Lc696              :in std_logic_vector(8 DOWNTO 0);
     Lc697              :in std_logic_vector(8 DOWNTO 0);
     Lc698              :in std_logic_vector(8 DOWNTO 0);
     Lc699              :in std_logic_vector(8 DOWNTO 0);
     Lc700              :in std_logic_vector(8 DOWNTO 0);
     Lc701              :in std_logic_vector(8 DOWNTO 0);
     Lc702              :in std_logic_vector(8 DOWNTO 0);
     Lc703              :in std_logic_vector(8 DOWNTO 0);
     Lc704              :in std_logic_vector(8 DOWNTO 0);
     Lc705              :in std_logic_vector(8 DOWNTO 0);
     Lc706              :in std_logic_vector(8 DOWNTO 0);
     Lc707              :in std_logic_vector(8 DOWNTO 0);
     Lc708              :in std_logic_vector(8 DOWNTO 0);
     Lc709              :in std_logic_vector(8 DOWNTO 0);
     Lc710              :in std_logic_vector(8 DOWNTO 0);
     Lc711              :in std_logic_vector(8 DOWNTO 0);
     Lc712              :in std_logic_vector(8 DOWNTO 0);
     Lc713              :in std_logic_vector(8 DOWNTO 0);
     Lc714              :in std_logic_vector(8 DOWNTO 0);
     Lc715              :in std_logic_vector(8 DOWNTO 0);
     Lc716              :in std_logic_vector(8 DOWNTO 0);
     Lc717              :in std_logic_vector(8 DOWNTO 0);
     Lc718              :in std_logic_vector(8 DOWNTO 0);
     Lc719              :in std_logic_vector(8 DOWNTO 0);
     Lc720              :in std_logic_vector(8 DOWNTO 0);
     Lc721              :in std_logic_vector(8 DOWNTO 0);
     Lc722              :in std_logic_vector(8 DOWNTO 0);
     Lc723              :in std_logic_vector(8 DOWNTO 0);
     Lc724              :in std_logic_vector(8 DOWNTO 0);
     Lc725              :in std_logic_vector(8 DOWNTO 0);
     Lc726              :in std_logic_vector(8 DOWNTO 0);
     Lc727              :in std_logic_vector(8 DOWNTO 0);
     Lc728              :in std_logic_vector(8 DOWNTO 0);
     Lc729              :in std_logic_vector(8 DOWNTO 0);
     Lc730              :in std_logic_vector(8 DOWNTO 0);
     Lc731              :in std_logic_vector(8 DOWNTO 0);
     Lc732              :in std_logic_vector(8 DOWNTO 0);
     Lc733              :in std_logic_vector(8 DOWNTO 0);
     Lc734              :in std_logic_vector(8 DOWNTO 0);
     Lc735              :in std_logic_vector(8 DOWNTO 0);
     Lc736              :in std_logic_vector(8 DOWNTO 0);
     Lc737              :in std_logic_vector(8 DOWNTO 0);
     Lc738              :in std_logic_vector(8 DOWNTO 0);
     Lc739              :in std_logic_vector(8 DOWNTO 0);
     Lc740              :in std_logic_vector(8 DOWNTO 0);
     Lc741              :in std_logic_vector(8 DOWNTO 0);
     Lc742              :in std_logic_vector(8 DOWNTO 0);
     Lc743              :in std_logic_vector(8 DOWNTO 0);
     Lc744              :in std_logic_vector(8 DOWNTO 0);
     Lc745              :in std_logic_vector(8 DOWNTO 0);
     Lc746              :in std_logic_vector(8 DOWNTO 0);
     Lc747              :in std_logic_vector(8 DOWNTO 0);
     Lc748              :in std_logic_vector(8 DOWNTO 0);
     Lc749              :in std_logic_vector(8 DOWNTO 0);
     Lc750              :in std_logic_vector(8 DOWNTO 0);
     Lc751              :in std_logic_vector(8 DOWNTO 0);
     Lc752              :in std_logic_vector(8 DOWNTO 0);
     Lc753              :in std_logic_vector(8 DOWNTO 0);
     Lc754              :in std_logic_vector(8 DOWNTO 0);
     Lc755              :in std_logic_vector(8 DOWNTO 0);
     Lc756              :in std_logic_vector(8 DOWNTO 0);
     Lc757              :in std_logic_vector(8 DOWNTO 0);
     Lc758              :in std_logic_vector(8 DOWNTO 0);
     Lc759              :in std_logic_vector(8 DOWNTO 0);
     Lc760              :in std_logic_vector(8 DOWNTO 0);
     Lc761              :in std_logic_vector(8 DOWNTO 0);
     Lc762              :in std_logic_vector(8 DOWNTO 0);
     Lc763              :in std_logic_vector(8 DOWNTO 0);
     Lc764              :in std_logic_vector(8 DOWNTO 0);
     Lc765              :in std_logic_vector(8 DOWNTO 0);
     Lc766              :in std_logic_vector(8 DOWNTO 0);
     Lc767              :in std_logic_vector(8 DOWNTO 0);
     Lc768              :in std_logic_vector(8 DOWNTO 0);
     Lc769              :in std_logic_vector(8 DOWNTO 0);
     Lc770              :in std_logic_vector(8 DOWNTO 0);
     Lc771              :in std_logic_vector(8 DOWNTO 0);
     Lc772              :in std_logic_vector(8 DOWNTO 0);
     Lc773              :in std_logic_vector(8 DOWNTO 0);
     Lc774              :in std_logic_vector(8 DOWNTO 0);
     Lc775              :in std_logic_vector(8 DOWNTO 0);
     Lc776              :in std_logic_vector(8 DOWNTO 0);
     Lc777              :in std_logic_vector(8 DOWNTO 0);
     Lc778              :in std_logic_vector(8 DOWNTO 0);
     Lc779              :in std_logic_vector(8 DOWNTO 0);
     Lc780              :in std_logic_vector(8 DOWNTO 0);
     Lc781              :in std_logic_vector(8 DOWNTO 0);
     Lc782              :in std_logic_vector(8 DOWNTO 0);
     Lc783              :in std_logic_vector(8 DOWNTO 0);
     Lc784              :in std_logic_vector(8 DOWNTO 0);
     Lc785              :in std_logic_vector(8 DOWNTO 0);
     Lc786              :in std_logic_vector(8 DOWNTO 0);
     Lc787              :in std_logic_vector(8 DOWNTO 0);
     Lc788              :in std_logic_vector(8 DOWNTO 0);
     Lc789              :in std_logic_vector(8 DOWNTO 0);
     Lc790              :in std_logic_vector(8 DOWNTO 0);
     Lc791              :in std_logic_vector(8 DOWNTO 0);
     Lc792              :in std_logic_vector(8 DOWNTO 0);
     Lc793              :in std_logic_vector(8 DOWNTO 0);
     Lc794              :in std_logic_vector(8 DOWNTO 0);
     Lc795              :in std_logic_vector(8 DOWNTO 0);
     Lc796              :in std_logic_vector(8 DOWNTO 0);
     Lc797              :in std_logic_vector(8 DOWNTO 0);
     Lc798              :in std_logic_vector(8 DOWNTO 0);
     Lc799              :in std_logic_vector(8 DOWNTO 0);
     Lc800              :in std_logic_vector(8 DOWNTO 0);
     Lc801              :in std_logic_vector(8 DOWNTO 0);
     Lc802              :in std_logic_vector(8 DOWNTO 0);
     Lc803              :in std_logic_vector(8 DOWNTO 0);
     Lc804              :in std_logic_vector(8 DOWNTO 0);
     Lc805              :in std_logic_vector(8 DOWNTO 0);
     Lc806              :in std_logic_vector(8 DOWNTO 0);
     Lc807              :in std_logic_vector(8 DOWNTO 0);
     Lc808              :in std_logic_vector(8 DOWNTO 0);
     Lc809              :in std_logic_vector(8 DOWNTO 0);
     Lc810              :in std_logic_vector(8 DOWNTO 0);
     Lc811              :in std_logic_vector(8 DOWNTO 0);
     Lc812              :in std_logic_vector(8 DOWNTO 0);
     Lc813              :in std_logic_vector(8 DOWNTO 0);
     Lc814              :in std_logic_vector(8 DOWNTO 0);
     Lc815              :in std_logic_vector(8 DOWNTO 0);
     Lc816              :in std_logic_vector(8 DOWNTO 0);
     Lc817              :in std_logic_vector(8 DOWNTO 0);
     Lc818              :in std_logic_vector(8 DOWNTO 0);
     Lc819              :in std_logic_vector(8 DOWNTO 0);
     Lc820              :in std_logic_vector(8 DOWNTO 0);
     Lc821              :in std_logic_vector(8 DOWNTO 0);
     Lc822              :in std_logic_vector(8 DOWNTO 0);
     Lc823              :in std_logic_vector(8 DOWNTO 0);
     Lc824              :in std_logic_vector(8 DOWNTO 0);
     Lc825              :in std_logic_vector(8 DOWNTO 0);
     Lc826              :in std_logic_vector(8 DOWNTO 0);
     Lc827              :in std_logic_vector(8 DOWNTO 0);
     Lc828              :in std_logic_vector(8 DOWNTO 0);
     Lc829              :in std_logic_vector(8 DOWNTO 0);
     Lc830              :in std_logic_vector(8 DOWNTO 0);
     Lc831              :in std_logic_vector(8 DOWNTO 0);
     Lc832              :in std_logic_vector(8 DOWNTO 0);
     Lc833              :in std_logic_vector(8 DOWNTO 0);
     Lc834              :in std_logic_vector(8 DOWNTO 0);
     Lc835              :in std_logic_vector(8 DOWNTO 0);
     Lc836              :in std_logic_vector(8 DOWNTO 0);
     Lc837              :in std_logic_vector(8 DOWNTO 0);
     Lc838              :in std_logic_vector(8 DOWNTO 0);
     Lc839              :in std_logic_vector(8 DOWNTO 0);
     Lc840              :in std_logic_vector(8 DOWNTO 0);
     Lc841              :in std_logic_vector(8 DOWNTO 0);
     Lc842              :in std_logic_vector(8 DOWNTO 0);
     Lc843              :in std_logic_vector(8 DOWNTO 0);
     Lc844              :in std_logic_vector(8 DOWNTO 0);
     Lc845              :in std_logic_vector(8 DOWNTO 0);
     Lc846              :in std_logic_vector(8 DOWNTO 0);
     Lc847              :in std_logic_vector(8 DOWNTO 0);
     Lc848              :in std_logic_vector(8 DOWNTO 0);
     Lc849              :in std_logic_vector(8 DOWNTO 0);
     Lc850              :in std_logic_vector(8 DOWNTO 0);
     Lc851              :in std_logic_vector(8 DOWNTO 0);
     Lc852              :in std_logic_vector(8 DOWNTO 0);
     Lc853              :in std_logic_vector(8 DOWNTO 0);
     Lc854              :in std_logic_vector(8 DOWNTO 0);
     Lc855              :in std_logic_vector(8 DOWNTO 0);
     Lc856              :in std_logic_vector(8 DOWNTO 0);
     Lc857              :in std_logic_vector(8 DOWNTO 0);
     Lc858              :in std_logic_vector(8 DOWNTO 0);
     Lc859              :in std_logic_vector(8 DOWNTO 0);
     Lc860              :in std_logic_vector(8 DOWNTO 0);
     Lc861              :in std_logic_vector(8 DOWNTO 0);
     Lc862              :in std_logic_vector(8 DOWNTO 0);
     Lc863              :in std_logic_vector(8 DOWNTO 0);
     Lc864              :in std_logic_vector(8 DOWNTO 0);
     Lc865              :in std_logic_vector(8 DOWNTO 0);
     Lc866              :in std_logic_vector(8 DOWNTO 0);
     Lc867              :in std_logic_vector(8 DOWNTO 0);
     Lc868              :in std_logic_vector(8 DOWNTO 0);
     Lc869              :in std_logic_vector(8 DOWNTO 0);
     Lc870              :in std_logic_vector(8 DOWNTO 0);
     Lc871              :in std_logic_vector(8 DOWNTO 0);
     Lc872              :in std_logic_vector(8 DOWNTO 0);
     Lc873              :in std_logic_vector(8 DOWNTO 0);
     Lc874              :in std_logic_vector(8 DOWNTO 0);
     Lc875              :in std_logic_vector(8 DOWNTO 0);
     Lc876              :in std_logic_vector(8 DOWNTO 0);
     Lc877              :in std_logic_vector(8 DOWNTO 0);
     Lc878              :in std_logic_vector(8 DOWNTO 0);
     Lc879              :in std_logic_vector(8 DOWNTO 0);
     Lc880              :in std_logic_vector(8 DOWNTO 0);
     Lc881              :in std_logic_vector(8 DOWNTO 0);
     Lc882              :in std_logic_vector(8 DOWNTO 0);
     Lc883              :in std_logic_vector(8 DOWNTO 0);
     Lc884              :in std_logic_vector(8 DOWNTO 0);
     Lc885              :in std_logic_vector(8 DOWNTO 0);
     Lc886              :in std_logic_vector(8 DOWNTO 0);
     Lc887              :in std_logic_vector(8 DOWNTO 0);
     Lc888              :in std_logic_vector(8 DOWNTO 0);
     Lc889              :in std_logic_vector(8 DOWNTO 0);
     Lc890              :in std_logic_vector(8 DOWNTO 0);
     Lc891              :in std_logic_vector(8 DOWNTO 0);
     Lc892              :in std_logic_vector(8 DOWNTO 0);
     Lc893              :in std_logic_vector(8 DOWNTO 0);
     Lc894              :in std_logic_vector(8 DOWNTO 0);
     Lc895              :in std_logic_vector(8 DOWNTO 0);
     Lc896              :in std_logic_vector(8 DOWNTO 0);
     Lc897              :in std_logic_vector(8 DOWNTO 0);
     Lc898              :in std_logic_vector(8 DOWNTO 0);
     Lc899              :in std_logic_vector(8 DOWNTO 0);
     Lc900              :in std_logic_vector(8 DOWNTO 0);
     Lc901              :in std_logic_vector(8 DOWNTO 0);
     Lc902              :in std_logic_vector(8 DOWNTO 0);
     Lc903              :in std_logic_vector(8 DOWNTO 0);
     Lc904              :in std_logic_vector(8 DOWNTO 0);
     Lc905              :in std_logic_vector(8 DOWNTO 0);
     Lc906              :in std_logic_vector(8 DOWNTO 0);
     Lc907              :in std_logic_vector(8 DOWNTO 0);
     Lc908              :in std_logic_vector(8 DOWNTO 0);
     Lc909              :in std_logic_vector(8 DOWNTO 0);
     Lc910              :in std_logic_vector(8 DOWNTO 0);
     Lc911              :in std_logic_vector(8 DOWNTO 0);
     Lc912              :in std_logic_vector(8 DOWNTO 0);
     Lc913              :in std_logic_vector(8 DOWNTO 0);
     Lc914              :in std_logic_vector(8 DOWNTO 0);
     Lc915              :in std_logic_vector(8 DOWNTO 0);
     Lc916              :in std_logic_vector(8 DOWNTO 0);
     Lc917              :in std_logic_vector(8 DOWNTO 0);
     Lc918              :in std_logic_vector(8 DOWNTO 0);
     Lc919              :in std_logic_vector(8 DOWNTO 0);
     Lc920              :in std_logic_vector(8 DOWNTO 0);
     Lc921              :in std_logic_vector(8 DOWNTO 0);
     Lc922              :in std_logic_vector(8 DOWNTO 0);
     Lc923              :in std_logic_vector(8 DOWNTO 0);
     Lc924              :in std_logic_vector(8 DOWNTO 0);
     Lc925              :in std_logic_vector(8 DOWNTO 0);
     Lc926              :in std_logic_vector(8 DOWNTO 0);
     Lc927              :in std_logic_vector(8 DOWNTO 0);
     Lc928              :in std_logic_vector(8 DOWNTO 0);
     Lc929              :in std_logic_vector(8 DOWNTO 0);
     Lc930              :in std_logic_vector(8 DOWNTO 0);
     Lc931              :in std_logic_vector(8 DOWNTO 0);
     Lc932              :in std_logic_vector(8 DOWNTO 0);
     Lc933              :in std_logic_vector(8 DOWNTO 0);
     Lc934              :in std_logic_vector(8 DOWNTO 0);
     Lc935              :in std_logic_vector(8 DOWNTO 0);
     Lc936              :in std_logic_vector(8 DOWNTO 0);
     Lc937              :in std_logic_vector(8 DOWNTO 0);
     Lc938              :in std_logic_vector(8 DOWNTO 0);
     Lc939              :in std_logic_vector(8 DOWNTO 0);
     Lc940              :in std_logic_vector(8 DOWNTO 0);
     Lc941              :in std_logic_vector(8 DOWNTO 0);
     Lc942              :in std_logic_vector(8 DOWNTO 0);
     Lc943              :in std_logic_vector(8 DOWNTO 0);
     Lc944              :in std_logic_vector(8 DOWNTO 0);
     Lc945              :in std_logic_vector(8 DOWNTO 0);
     Lc946              :in std_logic_vector(8 DOWNTO 0);
     Lc947              :in std_logic_vector(8 DOWNTO 0);
     Lc948              :in std_logic_vector(8 DOWNTO 0);
     Lc949              :in std_logic_vector(8 DOWNTO 0);
     Lc950              :in std_logic_vector(8 DOWNTO 0);
     Lc951              :in std_logic_vector(8 DOWNTO 0);
     Lc952              :in std_logic_vector(8 DOWNTO 0);
     Lc953              :in std_logic_vector(8 DOWNTO 0);
     Lc954              :in std_logic_vector(8 DOWNTO 0);
     Lc955              :in std_logic_vector(8 DOWNTO 0);
     Lc956              :in std_logic_vector(8 DOWNTO 0);
     Lc957              :in std_logic_vector(8 DOWNTO 0);
     Lc958              :in std_logic_vector(8 DOWNTO 0);
     Lc959              :in std_logic_vector(8 DOWNTO 0);
     Lc960              :in std_logic_vector(8 DOWNTO 0);
     Lc961              :in std_logic_vector(8 DOWNTO 0);
     Lc962              :in std_logic_vector(8 DOWNTO 0);
     Lc963              :in std_logic_vector(8 DOWNTO 0);
     Lc964              :in std_logic_vector(8 DOWNTO 0);
     Lc965              :in std_logic_vector(8 DOWNTO 0);
     Lc966              :in std_logic_vector(8 DOWNTO 0);
     Lc967              :in std_logic_vector(8 DOWNTO 0);
     Lc968              :in std_logic_vector(8 DOWNTO 0);
     Lc969              :in std_logic_vector(8 DOWNTO 0);
     Lc970              :in std_logic_vector(8 DOWNTO 0);
     Lc971              :in std_logic_vector(8 DOWNTO 0);
     Lc972              :in std_logic_vector(8 DOWNTO 0);
     Lc973              :in std_logic_vector(8 DOWNTO 0);
     Lc974              :in std_logic_vector(8 DOWNTO 0);
     Lc975              :in std_logic_vector(8 DOWNTO 0);
     Lc976              :in std_logic_vector(8 DOWNTO 0);
     Lc977              :in std_logic_vector(8 DOWNTO 0);
     Lc978              :in std_logic_vector(8 DOWNTO 0);
     Lc979              :in std_logic_vector(8 DOWNTO 0);
     Lc980              :in std_logic_vector(8 DOWNTO 0);
     Lc981              :in std_logic_vector(8 DOWNTO 0);
     Lc982              :in std_logic_vector(8 DOWNTO 0);
     Lc983              :in std_logic_vector(8 DOWNTO 0);
     Lc984              :in std_logic_vector(8 DOWNTO 0);
     Lc985              :in std_logic_vector(8 DOWNTO 0);
     Lc986              :in std_logic_vector(8 DOWNTO 0);
     Lc987              :in std_logic_vector(8 DOWNTO 0);
     Lc988              :in std_logic_vector(8 DOWNTO 0);
     Lc989              :in std_logic_vector(8 DOWNTO 0);
     Lc990              :in std_logic_vector(8 DOWNTO 0);
     Lc991              :in std_logic_vector(8 DOWNTO 0);
     Lc992              :in std_logic_vector(8 DOWNTO 0);
     Lc993              :in std_logic_vector(8 DOWNTO 0);
     Lc994              :in std_logic_vector(8 DOWNTO 0);
     Lc995              :in std_logic_vector(8 DOWNTO 0);
     Lc996              :in std_logic_vector(8 DOWNTO 0);
     Lc997              :in std_logic_vector(8 DOWNTO 0);
     Lc998              :in std_logic_vector(8 DOWNTO 0);
     Lc999              :in std_logic_vector(8 DOWNTO 0);
     Lc1000              :in std_logic_vector(8 DOWNTO 0);
     Lc1001              :in std_logic_vector(8 DOWNTO 0);
     Lc1002              :in std_logic_vector(8 DOWNTO 0);
     Lc1003              :in std_logic_vector(8 DOWNTO 0);
     Lc1004              :in std_logic_vector(8 DOWNTO 0);
     Lc1005              :in std_logic_vector(8 DOWNTO 0);
     Lc1006              :in std_logic_vector(8 DOWNTO 0);
     Lc1007              :in std_logic_vector(8 DOWNTO 0);
     Lc1008              :in std_logic_vector(8 DOWNTO 0);
     Lc1009              :in std_logic_vector(8 DOWNTO 0);
     Lc1010              :in std_logic_vector(8 DOWNTO 0);
     Lc1011              :in std_logic_vector(8 DOWNTO 0);
     Lc1012              :in std_logic_vector(8 DOWNTO 0);
     Lc1013              :in std_logic_vector(8 DOWNTO 0);
     Lc1014              :in std_logic_vector(8 DOWNTO 0);
     Lc1015              :in std_logic_vector(8 DOWNTO 0);
     Lc1016              :in std_logic_vector(8 DOWNTO 0);
     Lc1017              :in std_logic_vector(8 DOWNTO 0);
     Lc1018              :in std_logic_vector(8 DOWNTO 0);
     Lc1019              :in std_logic_vector(8 DOWNTO 0);
     Lc1020              :in std_logic_vector(8 DOWNTO 0);
     Lc1021              :in std_logic_vector(8 DOWNTO 0);
     Lc1022              :in std_logic_vector(8 DOWNTO 0);
     Lc1023              :in std_logic_vector(8 DOWNTO 0);
     Lc1024              :in std_logic_vector(8 DOWNTO 0);
     Lc1025              :in std_logic_vector(8 DOWNTO 0);
     Lc1026              :in std_logic_vector(8 DOWNTO 0);
     Lc1027              :in std_logic_vector(8 DOWNTO 0);
     Lc1028              :in std_logic_vector(8 DOWNTO 0);
     Lc1029              :in std_logic_vector(8 DOWNTO 0);
     Lc1030              :in std_logic_vector(8 DOWNTO 0);
     Lc1031              :in std_logic_vector(8 DOWNTO 0);
     Lc1032              :in std_logic_vector(8 DOWNTO 0);
     Lc1033              :in std_logic_vector(8 DOWNTO 0);
     Lc1034              :in std_logic_vector(8 DOWNTO 0);
     Lc1035              :in std_logic_vector(8 DOWNTO 0);
     Lc1036              :in std_logic_vector(8 DOWNTO 0);
     Lc1037              :in std_logic_vector(8 DOWNTO 0);
     Lc1038              :in std_logic_vector(8 DOWNTO 0);
     Lc1039              :in std_logic_vector(8 DOWNTO 0);
     Lc1040              :in std_logic_vector(8 DOWNTO 0);
     Lc1041              :in std_logic_vector(8 DOWNTO 0);
     Lc1042              :in std_logic_vector(8 DOWNTO 0);
     Lc1043              :in std_logic_vector(8 DOWNTO 0);
     Lc1044              :in std_logic_vector(8 DOWNTO 0);
     Lc1045              :in std_logic_vector(8 DOWNTO 0);
     Lc1046              :in std_logic_vector(8 DOWNTO 0);
     Lc1047              :in std_logic_vector(8 DOWNTO 0);
     Lc1048              :in std_logic_vector(8 DOWNTO 0);
     Lc1049              :in std_logic_vector(8 DOWNTO 0);
     Lc1050              :in std_logic_vector(8 DOWNTO 0);
     Lc1051              :in std_logic_vector(8 DOWNTO 0);
     Lc1052              :in std_logic_vector(8 DOWNTO 0);
     Lc1053              :in std_logic_vector(8 DOWNTO 0);
     Lc1054              :in std_logic_vector(8 DOWNTO 0);
     Lc1055              :in std_logic_vector(8 DOWNTO 0);
     Lc1056              :in std_logic_vector(8 DOWNTO 0);
     Lc1057              :in std_logic_vector(8 DOWNTO 0);
     Lc1058              :in std_logic_vector(8 DOWNTO 0);
     Lc1059              :in std_logic_vector(8 DOWNTO 0);
     Lc1060              :in std_logic_vector(8 DOWNTO 0);
     Lc1061              :in std_logic_vector(8 DOWNTO 0);
     Lc1062              :in std_logic_vector(8 DOWNTO 0);
     Lc1063              :in std_logic_vector(8 DOWNTO 0);
     Lc1064              :in std_logic_vector(8 DOWNTO 0);
     Lc1065              :in std_logic_vector(8 DOWNTO 0);
     Lc1066              :in std_logic_vector(8 DOWNTO 0);
     Lc1067              :in std_logic_vector(8 DOWNTO 0);
     Lc1068              :in std_logic_vector(8 DOWNTO 0);
     Lc1069              :in std_logic_vector(8 DOWNTO 0);
     Lc1070              :in std_logic_vector(8 DOWNTO 0);
     Lc1071              :in std_logic_vector(8 DOWNTO 0);
     Lc1072              :in std_logic_vector(8 DOWNTO 0);
     Lc1073              :in std_logic_vector(8 DOWNTO 0);
     Lc1074              :in std_logic_vector(8 DOWNTO 0);
     Lc1075              :in std_logic_vector(8 DOWNTO 0);
     Lc1076              :in std_logic_vector(8 DOWNTO 0);
     Lc1077              :in std_logic_vector(8 DOWNTO 0);
     Lc1078              :in std_logic_vector(8 DOWNTO 0);
     Lc1079              :in std_logic_vector(8 DOWNTO 0);
     Lc1080              :in std_logic_vector(8 DOWNTO 0);
     Lc1081              :in std_logic_vector(8 DOWNTO 0);
     Lc1082              :in std_logic_vector(8 DOWNTO 0);
     Lc1083              :in std_logic_vector(8 DOWNTO 0);
     Lc1084              :in std_logic_vector(8 DOWNTO 0);
     Lc1085              :in std_logic_vector(8 DOWNTO 0);
     Lc1086              :in std_logic_vector(8 DOWNTO 0);
     Lc1087              :in std_logic_vector(8 DOWNTO 0);
     Lc1088              :in std_logic_vector(8 DOWNTO 0);
     Lc1089              :in std_logic_vector(8 DOWNTO 0);
     Lc1090              :in std_logic_vector(8 DOWNTO 0);
     Lc1091              :in std_logic_vector(8 DOWNTO 0);
     Lc1092              :in std_logic_vector(8 DOWNTO 0);
     Lc1093              :in std_logic_vector(8 DOWNTO 0);
     Lc1094              :in std_logic_vector(8 DOWNTO 0);
     Lc1095              :in std_logic_vector(8 DOWNTO 0);
     Lc1096              :in std_logic_vector(8 DOWNTO 0);
     Lc1097              :in std_logic_vector(8 DOWNTO 0);
     Lc1098              :in std_logic_vector(8 DOWNTO 0);
     Lc1099              :in std_logic_vector(8 DOWNTO 0);
     Lc1100              :in std_logic_vector(8 DOWNTO 0);
     Lc1101              :in std_logic_vector(8 DOWNTO 0);
     Lc1102              :in std_logic_vector(8 DOWNTO 0);
     Lc1103              :in std_logic_vector(8 DOWNTO 0);
     Lc1104              :in std_logic_vector(8 DOWNTO 0);
     Lc1105              :in std_logic_vector(8 DOWNTO 0);
     Lc1106              :in std_logic_vector(8 DOWNTO 0);
     Lc1107              :in std_logic_vector(8 DOWNTO 0);
     Lc1108              :in std_logic_vector(8 DOWNTO 0);
     Lc1109              :in std_logic_vector(8 DOWNTO 0);
     Lc1110              :in std_logic_vector(8 DOWNTO 0);
     Lc1111              :in std_logic_vector(8 DOWNTO 0);
     Lc1112              :in std_logic_vector(8 DOWNTO 0);
     Lc1113              :in std_logic_vector(8 DOWNTO 0);
     Lc1114              :in std_logic_vector(8 DOWNTO 0);
     Lc1115              :in std_logic_vector(8 DOWNTO 0);
     Lc1116              :in std_logic_vector(8 DOWNTO 0);
     Lc1117              :in std_logic_vector(8 DOWNTO 0);
     Lc1118              :in std_logic_vector(8 DOWNTO 0);
     Lc1119              :in std_logic_vector(8 DOWNTO 0);
     Lc1120              :in std_logic_vector(8 DOWNTO 0);
     Lc1121              :in std_logic_vector(8 DOWNTO 0);
     Lc1122              :in std_logic_vector(8 DOWNTO 0);
     Lc1123              :in std_logic_vector(8 DOWNTO 0);
     Lc1124              :in std_logic_vector(8 DOWNTO 0);
     Lc1125              :in std_logic_vector(8 DOWNTO 0);
     Lc1126              :in std_logic_vector(8 DOWNTO 0);
     Lc1127              :in std_logic_vector(8 DOWNTO 0);
     Lc1128              :in std_logic_vector(8 DOWNTO 0);
     Lc1129              :in std_logic_vector(8 DOWNTO 0);
     Lc1130              :in std_logic_vector(8 DOWNTO 0);
     Lc1131              :in std_logic_vector(8 DOWNTO 0);
     Lc1132              :in std_logic_vector(8 DOWNTO 0);
     Lc1133              :in std_logic_vector(8 DOWNTO 0);
     Lc1134              :in std_logic_vector(8 DOWNTO 0);
     Lc1135              :in std_logic_vector(8 DOWNTO 0);
     Lc1136              :in std_logic_vector(8 DOWNTO 0);
     Lc1137              :in std_logic_vector(8 DOWNTO 0);
     Lc1138              :in std_logic_vector(8 DOWNTO 0);
     Lc1139              :in std_logic_vector(8 DOWNTO 0);
     Lc1140              :in std_logic_vector(8 DOWNTO 0);
     Lc1141              :in std_logic_vector(8 DOWNTO 0);
     Lc1142              :in std_logic_vector(8 DOWNTO 0);
     Lc1143              :in std_logic_vector(8 DOWNTO 0);
     Lc1144              :in std_logic_vector(8 DOWNTO 0);
     Lc1145              :in std_logic_vector(8 DOWNTO 0);
     Lc1146              :in std_logic_vector(8 DOWNTO 0);
     Lc1147              :in std_logic_vector(8 DOWNTO 0);
     Lc1148              :in std_logic_vector(8 DOWNTO 0);
     Lc1149              :in std_logic_vector(8 DOWNTO 0);
     Lc1150              :in std_logic_vector(8 DOWNTO 0);
     Lc1151              :in std_logic_vector(8 DOWNTO 0);
     Lc1152              :in std_logic_vector(8 DOWNTO 0);
     Lc1153              :in std_logic_vector(8 DOWNTO 0);
     Lc1154              :in std_logic_vector(8 DOWNTO 0);
     Lc1155              :in std_logic_vector(8 DOWNTO 0);
     Lc1156              :in std_logic_vector(8 DOWNTO 0);
     Lc1157              :in std_logic_vector(8 DOWNTO 0);
     Lc1158              :in std_logic_vector(8 DOWNTO 0);
     Lc1159              :in std_logic_vector(8 DOWNTO 0);
     Lc1160              :in std_logic_vector(8 DOWNTO 0);
     Lc1161              :in std_logic_vector(8 DOWNTO 0);
     Lc1162              :in std_logic_vector(8 DOWNTO 0);
     Lc1163              :in std_logic_vector(8 DOWNTO 0);
     Lc1164              :in std_logic_vector(8 DOWNTO 0);
     Lc1165              :in std_logic_vector(8 DOWNTO 0);
     Lc1166              :in std_logic_vector(8 DOWNTO 0);
     Lc1167              :in std_logic_vector(8 DOWNTO 0);
     Lc1168              :in std_logic_vector(8 DOWNTO 0);
     Lc1169              :in std_logic_vector(8 DOWNTO 0);
     Lc1170              :in std_logic_vector(8 DOWNTO 0);
     Lc1171              :in std_logic_vector(8 DOWNTO 0);
     Lc1172              :in std_logic_vector(8 DOWNTO 0);
     Lc1173              :in std_logic_vector(8 DOWNTO 0);
     Lc1174              :in std_logic_vector(8 DOWNTO 0);
     Lc1175              :in std_logic_vector(8 DOWNTO 0);
     Lc1176              :in std_logic_vector(8 DOWNTO 0);
     Lc1177              :in std_logic_vector(8 DOWNTO 0);
     Lc1178              :in std_logic_vector(8 DOWNTO 0);
     Lc1179              :in std_logic_vector(8 DOWNTO 0);
     Lc1180              :in std_logic_vector(8 DOWNTO 0);
     Lc1181              :in std_logic_vector(8 DOWNTO 0);
     Lc1182              :in std_logic_vector(8 DOWNTO 0);
     Lc1183              :in std_logic_vector(8 DOWNTO 0);
     Lc1184              :in std_logic_vector(8 DOWNTO 0);
     Lc1185              :in std_logic_vector(8 DOWNTO 0);
     Lc1186              :in std_logic_vector(8 DOWNTO 0);
     Lc1187              :in std_logic_vector(8 DOWNTO 0);
     Lc1188              :in std_logic_vector(8 DOWNTO 0);
     Lc1189              :in std_logic_vector(8 DOWNTO 0);
     Lc1190              :in std_logic_vector(8 DOWNTO 0);
     Lc1191              :in std_logic_vector(8 DOWNTO 0);
     Lc1192              :in std_logic_vector(8 DOWNTO 0);
     Lc1193              :in std_logic_vector(8 DOWNTO 0);
     Lc1194              :in std_logic_vector(8 DOWNTO 0);
     Lc1195              :in std_logic_vector(8 DOWNTO 0);
     Lc1196              :in std_logic_vector(8 DOWNTO 0);
     Lc1197              :in std_logic_vector(8 DOWNTO 0);
     Lc1198              :in std_logic_vector(8 DOWNTO 0);
     Lc1199              :in std_logic_vector(8 DOWNTO 0);
     Lc1200              :in std_logic_vector(8 DOWNTO 0);
     Lc1201              :in std_logic_vector(8 DOWNTO 0);
     Lc1202              :in std_logic_vector(8 DOWNTO 0);
     Lc1203              :in std_logic_vector(8 DOWNTO 0);
     Lc1204              :in std_logic_vector(8 DOWNTO 0);
     Lc1205              :in std_logic_vector(8 DOWNTO 0);
     Lc1206              :in std_logic_vector(8 DOWNTO 0);
     Lc1207              :in std_logic_vector(8 DOWNTO 0);
     Lc1208              :in std_logic_vector(8 DOWNTO 0);
     Lc1209              :in std_logic_vector(8 DOWNTO 0);
     Lc1210              :in std_logic_vector(8 DOWNTO 0);
     Lc1211              :in std_logic_vector(8 DOWNTO 0);
     Lc1212              :in std_logic_vector(8 DOWNTO 0);
     Lc1213              :in std_logic_vector(8 DOWNTO 0);
     Lc1214              :in std_logic_vector(8 DOWNTO 0);
     Lc1215              :in std_logic_vector(8 DOWNTO 0);
     Lc1216              :in std_logic_vector(8 DOWNTO 0);
     Lc1217              :in std_logic_vector(8 DOWNTO 0);
     Lc1218              :in std_logic_vector(8 DOWNTO 0);
     Lc1219              :in std_logic_vector(8 DOWNTO 0);
     Lc1220              :in std_logic_vector(8 DOWNTO 0);
     Lc1221              :in std_logic_vector(8 DOWNTO 0);
     Lc1222              :in std_logic_vector(8 DOWNTO 0);
     Lc1223              :in std_logic_vector(8 DOWNTO 0);
     Lc1224              :in std_logic_vector(8 DOWNTO 0);
     Lc1225              :in std_logic_vector(8 DOWNTO 0);
     Lc1226              :in std_logic_vector(8 DOWNTO 0);
     Lc1227              :in std_logic_vector(8 DOWNTO 0);
     Lc1228              :in std_logic_vector(8 DOWNTO 0);
     Lc1229              :in std_logic_vector(8 DOWNTO 0);
     Lc1230              :in std_logic_vector(8 DOWNTO 0);
     Lc1231              :in std_logic_vector(8 DOWNTO 0);
     Lc1232              :in std_logic_vector(8 DOWNTO 0);
     Lc1233              :in std_logic_vector(8 DOWNTO 0);
     Lc1234              :in std_logic_vector(8 DOWNTO 0);
     Lc1235              :in std_logic_vector(8 DOWNTO 0);
     Lc1236              :in std_logic_vector(8 DOWNTO 0);
     Lc1237              :in std_logic_vector(8 DOWNTO 0);
     Lc1238              :in std_logic_vector(8 DOWNTO 0);
     Lc1239              :in std_logic_vector(8 DOWNTO 0);
     Lc1240              :in std_logic_vector(8 DOWNTO 0);
     Lc1241              :in std_logic_vector(8 DOWNTO 0);
     Lc1242              :in std_logic_vector(8 DOWNTO 0);
     Lc1243              :in std_logic_vector(8 DOWNTO 0);
     Lc1244              :in std_logic_vector(8 DOWNTO 0);
     Lc1245              :in std_logic_vector(8 DOWNTO 0);
     Lc1246              :in std_logic_vector(8 DOWNTO 0);
     Lc1247              :in std_logic_vector(8 DOWNTO 0);
     Lc1248              :in std_logic_vector(8 DOWNTO 0);
     Lc1249              :in std_logic_vector(8 DOWNTO 0);
     Lc1250              :in std_logic_vector(8 DOWNTO 0);
     Lc1251              :in std_logic_vector(8 DOWNTO 0);
     Lc1252              :in std_logic_vector(8 DOWNTO 0);
     Lc1253              :in std_logic_vector(8 DOWNTO 0);
     Lc1254              :in std_logic_vector(8 DOWNTO 0);
     Lc1255              :in std_logic_vector(8 DOWNTO 0);
     Lc1256              :in std_logic_vector(8 DOWNTO 0);
     Lc1257              :in std_logic_vector(8 DOWNTO 0);
     Lc1258              :in std_logic_vector(8 DOWNTO 0);
     Lc1259              :in std_logic_vector(8 DOWNTO 0);
     Lc1260              :in std_logic_vector(8 DOWNTO 0);
     Lc1261              :in std_logic_vector(8 DOWNTO 0);
     Lc1262              :in std_logic_vector(8 DOWNTO 0);
     Lc1263              :in std_logic_vector(8 DOWNTO 0);
     Lc1264              :in std_logic_vector(8 DOWNTO 0);
     Lc1265              :in std_logic_vector(8 DOWNTO 0);
     Lc1266              :in std_logic_vector(8 DOWNTO 0);
     Lc1267              :in std_logic_vector(8 DOWNTO 0);
     Lc1268              :in std_logic_vector(8 DOWNTO 0);
     Lc1269              :in std_logic_vector(8 DOWNTO 0);
     Lc1270              :in std_logic_vector(8 DOWNTO 0);
     Lc1271              :in std_logic_vector(8 DOWNTO 0);
     Lc1272              :in std_logic_vector(8 DOWNTO 0);
     Lc1273              :in std_logic_vector(8 DOWNTO 0);
     Lc1274              :in std_logic_vector(8 DOWNTO 0);
     Lc1275              :in std_logic_vector(8 DOWNTO 0);
     Lc1276              :in std_logic_vector(8 DOWNTO 0);
     Lc1277              :in std_logic_vector(8 DOWNTO 0);
     Lc1278              :in std_logic_vector(8 DOWNTO 0);
     Lc1279              :in std_logic_vector(8 DOWNTO 0);
     Lc1280              :in std_logic_vector(8 DOWNTO 0);
     Lc1281              :in std_logic_vector(8 DOWNTO 0);
     Lc1282              :in std_logic_vector(8 DOWNTO 0);
     Lc1283              :in std_logic_vector(8 DOWNTO 0);
     Lc1284              :in std_logic_vector(8 DOWNTO 0);
     Lc1285              :in std_logic_vector(8 DOWNTO 0);
     Lc1286              :in std_logic_vector(8 DOWNTO 0);
     Lc1287              :in std_logic_vector(8 DOWNTO 0);
     Lc1288              :in std_logic_vector(8 DOWNTO 0);
     Lc1289              :in std_logic_vector(8 DOWNTO 0);
     Lc1290              :in std_logic_vector(8 DOWNTO 0);
     Lc1291              :in std_logic_vector(8 DOWNTO 0);
     Lc1292              :in std_logic_vector(8 DOWNTO 0);
     Lc1293              :in std_logic_vector(8 DOWNTO 0);
     Lc1294              :in std_logic_vector(8 DOWNTO 0);
     Lc1295              :in std_logic_vector(8 DOWNTO 0);
     Lc1296              :in std_logic_vector(8 DOWNTO 0);
     Lc1297              :in std_logic_vector(8 DOWNTO 0);
     Lc1298              :in std_logic_vector(8 DOWNTO 0);
     Lc1299              :in std_logic_vector(8 DOWNTO 0);
     Lc1300              :in std_logic_vector(8 DOWNTO 0);
     Lc1301              :in std_logic_vector(8 DOWNTO 0);
     Lc1302              :in std_logic_vector(8 DOWNTO 0);
     Lc1303              :in std_logic_vector(8 DOWNTO 0);
     Lc1304              :in std_logic_vector(8 DOWNTO 0);
     Lc1305              :in std_logic_vector(8 DOWNTO 0);
     Lc1306              :in std_logic_vector(8 DOWNTO 0);
     Lc1307              :in std_logic_vector(8 DOWNTO 0);
     Lc1308              :in std_logic_vector(8 DOWNTO 0);
     Lc1309              :in std_logic_vector(8 DOWNTO 0);
     Lc1310              :in std_logic_vector(8 DOWNTO 0);
     Lc1311              :in std_logic_vector(8 DOWNTO 0);
     Lc1312              :in std_logic_vector(8 DOWNTO 0);
     Lc1313              :in std_logic_vector(8 DOWNTO 0);
     Lc1314              :in std_logic_vector(8 DOWNTO 0);
     Lc1315              :in std_logic_vector(8 DOWNTO 0);
     Lc1316              :in std_logic_vector(8 DOWNTO 0);
     Lc1317              :in std_logic_vector(8 DOWNTO 0);
     Lc1318              :in std_logic_vector(8 DOWNTO 0);
     Lc1319              :in std_logic_vector(8 DOWNTO 0);
     Lc1320              :in std_logic_vector(8 DOWNTO 0);
     Lc1321              :in std_logic_vector(8 DOWNTO 0);
     Lc1322              :in std_logic_vector(8 DOWNTO 0);
     Lc1323              :in std_logic_vector(8 DOWNTO 0);
     Lc1324              :in std_logic_vector(8 DOWNTO 0);
     Lc1325              :in std_logic_vector(8 DOWNTO 0);
     Lc1326              :in std_logic_vector(8 DOWNTO 0);
     Lc1327              :in std_logic_vector(8 DOWNTO 0);
     Lc1328              :in std_logic_vector(8 DOWNTO 0);
     Lc1329              :in std_logic_vector(8 DOWNTO 0);
     Lc1330              :in std_logic_vector(8 DOWNTO 0);
     Lc1331              :in std_logic_vector(8 DOWNTO 0);
     Lc1332              :in std_logic_vector(8 DOWNTO 0);
     Lc1333              :in std_logic_vector(8 DOWNTO 0);
     Lc1334              :in std_logic_vector(8 DOWNTO 0);
     Lc1335              :in std_logic_vector(8 DOWNTO 0);
     Lc1336              :in std_logic_vector(8 DOWNTO 0);
     Lc1337              :in std_logic_vector(8 DOWNTO 0);
     Lc1338              :in std_logic_vector(8 DOWNTO 0);
     Lc1339              :in std_logic_vector(8 DOWNTO 0);
     Lc1340              :in std_logic_vector(8 DOWNTO 0);
     Lc1341              :in std_logic_vector(8 DOWNTO 0);
     Lc1342              :in std_logic_vector(8 DOWNTO 0);
     Lc1343              :in std_logic_vector(8 DOWNTO 0);
     Lc1344              :in std_logic_vector(8 DOWNTO 0);
     Lc1345              :in std_logic_vector(8 DOWNTO 0);
     Lc1346              :in std_logic_vector(8 DOWNTO 0);
     Lc1347              :in std_logic_vector(8 DOWNTO 0);
     Lc1348              :in std_logic_vector(8 DOWNTO 0);
     Lc1349              :in std_logic_vector(8 DOWNTO 0);
     Lc1350              :in std_logic_vector(8 DOWNTO 0);
     Lc1351              :in std_logic_vector(8 DOWNTO 0);
     Lc1352              :in std_logic_vector(8 DOWNTO 0);
     Lc1353              :in std_logic_vector(8 DOWNTO 0);
     Lc1354              :in std_logic_vector(8 DOWNTO 0);
     Lc1355              :in std_logic_vector(8 DOWNTO 0);
     Lc1356              :in std_logic_vector(8 DOWNTO 0);
     Lc1357              :in std_logic_vector(8 DOWNTO 0);
     Lc1358              :in std_logic_vector(8 DOWNTO 0);
     Lc1359              :in std_logic_vector(8 DOWNTO 0);
     Lc1360              :in std_logic_vector(8 DOWNTO 0);
     Lc1361              :in std_logic_vector(8 DOWNTO 0);
     Lc1362              :in std_logic_vector(8 DOWNTO 0);
     Lc1363              :in std_logic_vector(8 DOWNTO 0);
     Lc1364              :in std_logic_vector(8 DOWNTO 0);
     Lc1365              :in std_logic_vector(8 DOWNTO 0);
     Lc1366              :in std_logic_vector(8 DOWNTO 0);
     Lc1367              :in std_logic_vector(8 DOWNTO 0);
     Lc1368              :in std_logic_vector(8 DOWNTO 0);
     Lc1369              :in std_logic_vector(8 DOWNTO 0);
     Lc1370              :in std_logic_vector(8 DOWNTO 0);
     Lc1371              :in std_logic_vector(8 DOWNTO 0);
     Lc1372              :in std_logic_vector(8 DOWNTO 0);
     Lc1373              :in std_logic_vector(8 DOWNTO 0);
     Lc1374              :in std_logic_vector(8 DOWNTO 0);
     Lc1375              :in std_logic_vector(8 DOWNTO 0);
     Lc1376              :in std_logic_vector(8 DOWNTO 0);
     Lc1377              :in std_logic_vector(8 DOWNTO 0);
     Lc1378              :in std_logic_vector(8 DOWNTO 0);
     Lc1379              :in std_logic_vector(8 DOWNTO 0);
     Lc1380              :in std_logic_vector(8 DOWNTO 0);
     Lc1381              :in std_logic_vector(8 DOWNTO 0);
     Lc1382              :in std_logic_vector(8 DOWNTO 0);
     Lc1383              :in std_logic_vector(8 DOWNTO 0);
     Lc1384              :in std_logic_vector(8 DOWNTO 0);
     Lc1385              :in std_logic_vector(8 DOWNTO 0);
     Lc1386              :in std_logic_vector(8 DOWNTO 0);
     Lc1387              :in std_logic_vector(8 DOWNTO 0);
     Lc1388              :in std_logic_vector(8 DOWNTO 0);
     Lc1389              :in std_logic_vector(8 DOWNTO 0);
     Lc1390              :in std_logic_vector(8 DOWNTO 0);
     Lc1391              :in std_logic_vector(8 DOWNTO 0);
     Lc1392              :in std_logic_vector(8 DOWNTO 0);
     Lc1393              :in std_logic_vector(8 DOWNTO 0);
     Lc1394              :in std_logic_vector(8 DOWNTO 0);
     Lc1395              :in std_logic_vector(8 DOWNTO 0);
     Lc1396              :in std_logic_vector(8 DOWNTO 0);
     Lc1397              :in std_logic_vector(8 DOWNTO 0);
     Lc1398              :in std_logic_vector(8 DOWNTO 0);
     Lc1399              :in std_logic_vector(8 DOWNTO 0);
     Lc1400              :in std_logic_vector(8 DOWNTO 0);
     Lc1401              :in std_logic_vector(8 DOWNTO 0);
     Lc1402              :in std_logic_vector(8 DOWNTO 0);
     Lc1403              :in std_logic_vector(8 DOWNTO 0);
     Lc1404              :in std_logic_vector(8 DOWNTO 0);
     Lc1405              :in std_logic_vector(8 DOWNTO 0);
     Lc1406              :in std_logic_vector(8 DOWNTO 0);
     Lc1407              :in std_logic_vector(8 DOWNTO 0);
     Lc1408              :in std_logic_vector(8 DOWNTO 0);
     Lc1409              :in std_logic_vector(8 DOWNTO 0);
     Lc1410              :in std_logic_vector(8 DOWNTO 0);
     Lc1411              :in std_logic_vector(8 DOWNTO 0);
     Lc1412              :in std_logic_vector(8 DOWNTO 0);
     Lc1413              :in std_logic_vector(8 DOWNTO 0);
     Lc1414              :in std_logic_vector(8 DOWNTO 0);
     Lc1415              :in std_logic_vector(8 DOWNTO 0);
     Lc1416              :in std_logic_vector(8 DOWNTO 0);
     Lc1417              :in std_logic_vector(8 DOWNTO 0);
     Lc1418              :in std_logic_vector(8 DOWNTO 0);
     Lc1419              :in std_logic_vector(8 DOWNTO 0);
     Lc1420              :in std_logic_vector(8 DOWNTO 0);
     Lc1421              :in std_logic_vector(8 DOWNTO 0);
     Lc1422              :in std_logic_vector(8 DOWNTO 0);
     Lc1423              :in std_logic_vector(8 DOWNTO 0);
     Lc1424              :in std_logic_vector(8 DOWNTO 0);
     Lc1425              :in std_logic_vector(8 DOWNTO 0);
     Lc1426              :in std_logic_vector(8 DOWNTO 0);
     Lc1427              :in std_logic_vector(8 DOWNTO 0);
     Lc1428              :in std_logic_vector(8 DOWNTO 0);
     Lc1429              :in std_logic_vector(8 DOWNTO 0);
     Lc1430              :in std_logic_vector(8 DOWNTO 0);
     Lc1431              :in std_logic_vector(8 DOWNTO 0);
     Lc1432              :in std_logic_vector(8 DOWNTO 0);
     Lc1433              :in std_logic_vector(8 DOWNTO 0);
     Lc1434              :in std_logic_vector(8 DOWNTO 0);
     Lc1435              :in std_logic_vector(8 DOWNTO 0);
     Lc1436              :in std_logic_vector(8 DOWNTO 0);
     Lc1437              :in std_logic_vector(8 DOWNTO 0);
     Lc1438              :in std_logic_vector(8 DOWNTO 0);
     Lc1439              :in std_logic_vector(8 DOWNTO 0);
     Lc1440              :in std_logic_vector(8 DOWNTO 0);
     Lc1441              :in std_logic_vector(8 DOWNTO 0);
     Lc1442              :in std_logic_vector(8 DOWNTO 0);
     Lc1443              :in std_logic_vector(8 DOWNTO 0);
     Lc1444              :in std_logic_vector(8 DOWNTO 0);
     Lc1445              :in std_logic_vector(8 DOWNTO 0);
     Lc1446              :in std_logic_vector(8 DOWNTO 0);
     Lc1447              :in std_logic_vector(8 DOWNTO 0);
     Lc1448              :in std_logic_vector(8 DOWNTO 0);
     Lc1449              :in std_logic_vector(8 DOWNTO 0);
     Lc1450              :in std_logic_vector(8 DOWNTO 0);
     Lc1451              :in std_logic_vector(8 DOWNTO 0);
     Lc1452              :in std_logic_vector(8 DOWNTO 0);
     Lc1453              :in std_logic_vector(8 DOWNTO 0);
     Lc1454              :in std_logic_vector(8 DOWNTO 0);
     Lc1455              :in std_logic_vector(8 DOWNTO 0);
     Lc1456              :in std_logic_vector(8 DOWNTO 0);
     Lc1457              :in std_logic_vector(8 DOWNTO 0);
     Lc1458              :in std_logic_vector(8 DOWNTO 0);
     Lc1459              :in std_logic_vector(8 DOWNTO 0);
     Lc1460              :in std_logic_vector(8 DOWNTO 0);
     Lc1461              :in std_logic_vector(8 DOWNTO 0);
     Lc1462              :in std_logic_vector(8 DOWNTO 0);
     Lc1463              :in std_logic_vector(8 DOWNTO 0);
     Lc1464              :in std_logic_vector(8 DOWNTO 0);
     Lc1465              :in std_logic_vector(8 DOWNTO 0);
     Lc1466              :in std_logic_vector(8 DOWNTO 0);
     Lc1467              :in std_logic_vector(8 DOWNTO 0);
     Lc1468              :in std_logic_vector(8 DOWNTO 0);
     Lc1469              :in std_logic_vector(8 DOWNTO 0);
     Lc1470              :in std_logic_vector(8 DOWNTO 0);
     Lc1471              :in std_logic_vector(8 DOWNTO 0);
     Lc1472              :in std_logic_vector(8 DOWNTO 0);
     Lc1473              :in std_logic_vector(8 DOWNTO 0);
     Lc1474              :in std_logic_vector(8 DOWNTO 0);
     Lc1475              :in std_logic_vector(8 DOWNTO 0);
     Lc1476              :in std_logic_vector(8 DOWNTO 0);
     Lc1477              :in std_logic_vector(8 DOWNTO 0);
     Lc1478              :in std_logic_vector(8 DOWNTO 0);
     Lc1479              :in std_logic_vector(8 DOWNTO 0);
     Lc1480              :in std_logic_vector(8 DOWNTO 0);
     Lc1481              :in std_logic_vector(8 DOWNTO 0);
     Lc1482              :in std_logic_vector(8 DOWNTO 0);
     Lc1483              :in std_logic_vector(8 DOWNTO 0);
     Lc1484              :in std_logic_vector(8 DOWNTO 0);
     Lc1485              :in std_logic_vector(8 DOWNTO 0);
     Lc1486              :in std_logic_vector(8 DOWNTO 0);
     Lc1487              :in std_logic_vector(8 DOWNTO 0);
     Lc1488              :in std_logic_vector(8 DOWNTO 0);
     Lc1489              :in std_logic_vector(8 DOWNTO 0);
     Lc1490              :in std_logic_vector(8 DOWNTO 0);
     Lc1491              :in std_logic_vector(8 DOWNTO 0);
     Lc1492              :in std_logic_vector(8 DOWNTO 0);
     Lc1493              :in std_logic_vector(8 DOWNTO 0);
     Lc1494              :in std_logic_vector(8 DOWNTO 0);
     Lc1495              :in std_logic_vector(8 DOWNTO 0);
     Lc1496              :in std_logic_vector(8 DOWNTO 0);
     Lc1497              :in std_logic_vector(8 DOWNTO 0);
     Lc1498              :in std_logic_vector(8 DOWNTO 0);
     Lc1499              :in std_logic_vector(8 DOWNTO 0);
     Lc1500              :in std_logic_vector(8 DOWNTO 0);
     Lc1501              :in std_logic_vector(8 DOWNTO 0);
     Lc1502              :in std_logic_vector(8 DOWNTO 0);
     Lc1503              :in std_logic_vector(8 DOWNTO 0);
     Lc1504              :in std_logic_vector(8 DOWNTO 0);
     Lc1505              :in std_logic_vector(8 DOWNTO 0);
     Lc1506              :in std_logic_vector(8 DOWNTO 0);
     Lc1507              :in std_logic_vector(8 DOWNTO 0);
     Lc1508              :in std_logic_vector(8 DOWNTO 0);
     Lc1509              :in std_logic_vector(8 DOWNTO 0);
     Lc1510              :in std_logic_vector(8 DOWNTO 0);
     Lc1511              :in std_logic_vector(8 DOWNTO 0);
     Lc1512              :in std_logic_vector(8 DOWNTO 0);
     Lc1513              :in std_logic_vector(8 DOWNTO 0);
     Lc1514              :in std_logic_vector(8 DOWNTO 0);
     Lc1515              :in std_logic_vector(8 DOWNTO 0);
     Lc1516              :in std_logic_vector(8 DOWNTO 0);
     Lc1517              :in std_logic_vector(8 DOWNTO 0);
     Lc1518              :in std_logic_vector(8 DOWNTO 0);
     Lc1519              :in std_logic_vector(8 DOWNTO 0);
     Lc1520              :in std_logic_vector(8 DOWNTO 0);
     Lc1521              :in std_logic_vector(8 DOWNTO 0);
     Lc1522              :in std_logic_vector(8 DOWNTO 0);
     Lc1523              :in std_logic_vector(8 DOWNTO 0);
     Lc1524              :in std_logic_vector(8 DOWNTO 0);
     Lc1525              :in std_logic_vector(8 DOWNTO 0);
     Lc1526              :in std_logic_vector(8 DOWNTO 0);
     Lc1527              :in std_logic_vector(8 DOWNTO 0);
     Lc1528              :in std_logic_vector(8 DOWNTO 0);
     Lc1529              :in std_logic_vector(8 DOWNTO 0);
     Lc1530              :in std_logic_vector(8 DOWNTO 0);
     Lc1531              :in std_logic_vector(8 DOWNTO 0);
     Lc1532              :in std_logic_vector(8 DOWNTO 0);
     Lc1533              :in std_logic_vector(8 DOWNTO 0);
     Lc1534              :in std_logic_vector(8 DOWNTO 0);
     Lc1535              :in std_logic_vector(8 DOWNTO 0);
     Lc1536              :in std_logic_vector(8 DOWNTO 0);
     Lc1537              :in std_logic_vector(8 DOWNTO 0);
     Lc1538              :in std_logic_vector(8 DOWNTO 0);
     Lc1539              :in std_logic_vector(8 DOWNTO 0);
     Lc1540              :in std_logic_vector(8 DOWNTO 0);
     Lc1541              :in std_logic_vector(8 DOWNTO 0);
     Lc1542              :in std_logic_vector(8 DOWNTO 0);
     Lc1543              :in std_logic_vector(8 DOWNTO 0);
     Lc1544              :in std_logic_vector(8 DOWNTO 0);
     Lc1545              :in std_logic_vector(8 DOWNTO 0);
     Lc1546              :in std_logic_vector(8 DOWNTO 0);
     Lc1547              :in std_logic_vector(8 DOWNTO 0);
     Lc1548              :in std_logic_vector(8 DOWNTO 0);
     Lc1549              :in std_logic_vector(8 DOWNTO 0);
     Lc1550              :in std_logic_vector(8 DOWNTO 0);
     Lc1551              :in std_logic_vector(8 DOWNTO 0);
     Lc1552              :in std_logic_vector(8 DOWNTO 0);
     Lc1553              :in std_logic_vector(8 DOWNTO 0);
     Lc1554              :in std_logic_vector(8 DOWNTO 0);
     Lc1555              :in std_logic_vector(8 DOWNTO 0);
     Lc1556              :in std_logic_vector(8 DOWNTO 0);
     Lc1557              :in std_logic_vector(8 DOWNTO 0);
     Lc1558              :in std_logic_vector(8 DOWNTO 0);
     Lc1559              :in std_logic_vector(8 DOWNTO 0);
     Lc1560              :in std_logic_vector(8 DOWNTO 0);
     Lc1561              :in std_logic_vector(8 DOWNTO 0);
     Lc1562              :in std_logic_vector(8 DOWNTO 0);
     Lc1563              :in std_logic_vector(8 DOWNTO 0);
     Lc1564              :in std_logic_vector(8 DOWNTO 0);
     Lc1565              :in std_logic_vector(8 DOWNTO 0);
     Lc1566              :in std_logic_vector(8 DOWNTO 0);
     Lc1567              :in std_logic_vector(8 DOWNTO 0);
     Lc1568              :in std_logic_vector(8 DOWNTO 0);
     Lc1569              :in std_logic_vector(8 DOWNTO 0);
     Lc1570              :in std_logic_vector(8 DOWNTO 0);
     Lc1571              :in std_logic_vector(8 DOWNTO 0);
     Lc1572              :in std_logic_vector(8 DOWNTO 0);
     Lc1573              :in std_logic_vector(8 DOWNTO 0);
     Lc1574              :in std_logic_vector(8 DOWNTO 0);
     Lc1575              :in std_logic_vector(8 DOWNTO 0);
     Lc1576              :in std_logic_vector(8 DOWNTO 0);
     Lc1577              :in std_logic_vector(8 DOWNTO 0);
     Lc1578              :in std_logic_vector(8 DOWNTO 0);
     Lc1579              :in std_logic_vector(8 DOWNTO 0);
     Lc1580              :in std_logic_vector(8 DOWNTO 0);
     Lc1581              :in std_logic_vector(8 DOWNTO 0);
     Lc1582              :in std_logic_vector(8 DOWNTO 0);
     Lc1583              :in std_logic_vector(8 DOWNTO 0);
     Lc1584              :in std_logic_vector(8 DOWNTO 0);
     Lc1585              :in std_logic_vector(8 DOWNTO 0);
     Lc1586              :in std_logic_vector(8 DOWNTO 0);
     Lc1587              :in std_logic_vector(8 DOWNTO 0);
     Lc1588              :in std_logic_vector(8 DOWNTO 0);
     Lc1589              :in std_logic_vector(8 DOWNTO 0);
     Lc1590              :in std_logic_vector(8 DOWNTO 0);
     Lc1591              :in std_logic_vector(8 DOWNTO 0);
     Lc1592              :in std_logic_vector(8 DOWNTO 0);
     Lc1593              :in std_logic_vector(8 DOWNTO 0);
     Lc1594              :in std_logic_vector(8 DOWNTO 0);
     Lc1595              :in std_logic_vector(8 DOWNTO 0);
     Lc1596              :in std_logic_vector(8 DOWNTO 0);
     Lc1597              :in std_logic_vector(8 DOWNTO 0);
     Lc1598              :in std_logic_vector(8 DOWNTO 0);
     Lc1599              :in std_logic_vector(8 DOWNTO 0);
     Lc1600              :in std_logic_vector(8 DOWNTO 0);
     Lc1601              :in std_logic_vector(8 DOWNTO 0);
     Lc1602              :in std_logic_vector(8 DOWNTO 0);
     Lc1603              :in std_logic_vector(8 DOWNTO 0);
     Lc1604              :in std_logic_vector(8 DOWNTO 0);
     Lc1605              :in std_logic_vector(8 DOWNTO 0);
     Lc1606              :in std_logic_vector(8 DOWNTO 0);
     Lc1607              :in std_logic_vector(8 DOWNTO 0);
     Lc1608              :in std_logic_vector(8 DOWNTO 0);
     Lc1609              :in std_logic_vector(8 DOWNTO 0);
     Lc1610              :in std_logic_vector(8 DOWNTO 0);
     Lc1611              :in std_logic_vector(8 DOWNTO 0);
     Lc1612              :in std_logic_vector(8 DOWNTO 0);
     Lc1613              :in std_logic_vector(8 DOWNTO 0);
     Lc1614              :in std_logic_vector(8 DOWNTO 0);
     Lc1615              :in std_logic_vector(8 DOWNTO 0);
     Lc1616              :in std_logic_vector(8 DOWNTO 0);
     Lc1617              :in std_logic_vector(8 DOWNTO 0);
     Lc1618              :in std_logic_vector(8 DOWNTO 0);
     Lc1619              :in std_logic_vector(8 DOWNTO 0);
     Lc1620              :in std_logic_vector(8 DOWNTO 0);
     Lc1621              :in std_logic_vector(8 DOWNTO 0);
     Lc1622              :in std_logic_vector(8 DOWNTO 0);
     Lc1623              :in std_logic_vector(8 DOWNTO 0);
     Lc1624              :in std_logic_vector(8 DOWNTO 0);
     Lc1625              :in std_logic_vector(8 DOWNTO 0);
     Lc1626              :in std_logic_vector(8 DOWNTO 0);
     Lc1627              :in std_logic_vector(8 DOWNTO 0);
     Lc1628              :in std_logic_vector(8 DOWNTO 0);
     Lc1629              :in std_logic_vector(8 DOWNTO 0);
     Lc1630              :in std_logic_vector(8 DOWNTO 0);
     Lc1631              :in std_logic_vector(8 DOWNTO 0);
     Lc1632              :in std_logic_vector(8 DOWNTO 0);
     Lc1633              :in std_logic_vector(8 DOWNTO 0);
     Lc1634              :in std_logic_vector(8 DOWNTO 0);
     Lc1635              :in std_logic_vector(8 DOWNTO 0);
     Lc1636              :in std_logic_vector(8 DOWNTO 0);
     Lc1637              :in std_logic_vector(8 DOWNTO 0);
     Lc1638              :in std_logic_vector(8 DOWNTO 0);
     Lc1639              :in std_logic_vector(8 DOWNTO 0);
     Lc1640              :in std_logic_vector(8 DOWNTO 0);
     Lc1641              :in std_logic_vector(8 DOWNTO 0);
     Lc1642              :in std_logic_vector(8 DOWNTO 0);
     Lc1643              :in std_logic_vector(8 DOWNTO 0);
     Lc1644              :in std_logic_vector(8 DOWNTO 0);
     Lc1645              :in std_logic_vector(8 DOWNTO 0);
     Lc1646              :in std_logic_vector(8 DOWNTO 0);
     Lc1647              :in std_logic_vector(8 DOWNTO 0);
     Lc1648              :in std_logic_vector(8 DOWNTO 0);
     Lc1649              :in std_logic_vector(8 DOWNTO 0);
     Lc1650              :in std_logic_vector(8 DOWNTO 0);
     Lc1651              :in std_logic_vector(8 DOWNTO 0);
     Lc1652              :in std_logic_vector(8 DOWNTO 0);
     Lc1653              :in std_logic_vector(8 DOWNTO 0);
     Lc1654              :in std_logic_vector(8 DOWNTO 0);
     Lc1655              :in std_logic_vector(8 DOWNTO 0);
     Lc1656              :in std_logic_vector(8 DOWNTO 0);
     Lc1657              :in std_logic_vector(8 DOWNTO 0);
     Lc1658              :in std_logic_vector(8 DOWNTO 0);
     Lc1659              :in std_logic_vector(8 DOWNTO 0);
     Lc1660              :in std_logic_vector(8 DOWNTO 0);
     Lc1661              :in std_logic_vector(8 DOWNTO 0);
     Lc1662              :in std_logic_vector(8 DOWNTO 0);
     Lc1663              :in std_logic_vector(8 DOWNTO 0);
     Lc1664              :in std_logic_vector(8 DOWNTO 0);
     Lc1665              :in std_logic_vector(8 DOWNTO 0);
     Lc1666              :in std_logic_vector(8 DOWNTO 0);
     Lc1667              :in std_logic_vector(8 DOWNTO 0);
     Lc1668              :in std_logic_vector(8 DOWNTO 0);
     Lc1669              :in std_logic_vector(8 DOWNTO 0);
     Lc1670              :in std_logic_vector(8 DOWNTO 0);
     Lc1671              :in std_logic_vector(8 DOWNTO 0);
     Lc1672              :in std_logic_vector(8 DOWNTO 0);
     Lc1673              :in std_logic_vector(8 DOWNTO 0);
     Lc1674              :in std_logic_vector(8 DOWNTO 0);
     Lc1675              :in std_logic_vector(8 DOWNTO 0);
     Lc1676              :in std_logic_vector(8 DOWNTO 0);
     Lc1677              :in std_logic_vector(8 DOWNTO 0);
     Lc1678              :in std_logic_vector(8 DOWNTO 0);
     Lc1679              :in std_logic_vector(8 DOWNTO 0);
     Lc1680              :in std_logic_vector(8 DOWNTO 0);
     Lc1681              :in std_logic_vector(8 DOWNTO 0);
     Lc1682              :in std_logic_vector(8 DOWNTO 0);
     Lc1683              :in std_logic_vector(8 DOWNTO 0);
     Lc1684              :in std_logic_vector(8 DOWNTO 0);
     Lc1685              :in std_logic_vector(8 DOWNTO 0);
     Lc1686              :in std_logic_vector(8 DOWNTO 0);
     Lc1687              :in std_logic_vector(8 DOWNTO 0);
     Lc1688              :in std_logic_vector(8 DOWNTO 0);
     Lc1689              :in std_logic_vector(8 DOWNTO 0);
     Lc1690              :in std_logic_vector(8 DOWNTO 0);
     Lc1691              :in std_logic_vector(8 DOWNTO 0);
     Lc1692              :in std_logic_vector(8 DOWNTO 0);
     Lc1693              :in std_logic_vector(8 DOWNTO 0);
     Lc1694              :in std_logic_vector(8 DOWNTO 0);
     Lc1695              :in std_logic_vector(8 DOWNTO 0);
     Lc1696              :in std_logic_vector(8 DOWNTO 0);
     Lc1697              :in std_logic_vector(8 DOWNTO 0);
     Lc1698              :in std_logic_vector(8 DOWNTO 0);
     Lc1699              :in std_logic_vector(8 DOWNTO 0);
     Lc1700              :in std_logic_vector(8 DOWNTO 0);
     Lc1701              :in std_logic_vector(8 DOWNTO 0);
     Lc1702              :in std_logic_vector(8 DOWNTO 0);
     Lc1703              :in std_logic_vector(8 DOWNTO 0);
     Lc1704              :in std_logic_vector(8 DOWNTO 0);
     Lc1705              :in std_logic_vector(8 DOWNTO 0);
     Lc1706              :in std_logic_vector(8 DOWNTO 0);
     Lc1707              :in std_logic_vector(8 DOWNTO 0);
     Lc1708              :in std_logic_vector(8 DOWNTO 0);
     Lc1709              :in std_logic_vector(8 DOWNTO 0);
     Lc1710              :in std_logic_vector(8 DOWNTO 0);
     Lc1711              :in std_logic_vector(8 DOWNTO 0);
     Lc1712              :in std_logic_vector(8 DOWNTO 0);
     Lc1713              :in std_logic_vector(8 DOWNTO 0);
     Lc1714              :in std_logic_vector(8 DOWNTO 0);
     Lc1715              :in std_logic_vector(8 DOWNTO 0);
     Lc1716              :in std_logic_vector(8 DOWNTO 0);
     Lc1717              :in std_logic_vector(8 DOWNTO 0);
     Lc1718              :in std_logic_vector(8 DOWNTO 0);
     Lc1719              :in std_logic_vector(8 DOWNTO 0);
     Lc1720              :in std_logic_vector(8 DOWNTO 0);
     Lc1721              :in std_logic_vector(8 DOWNTO 0);
     Lc1722              :in std_logic_vector(8 DOWNTO 0);
     Lc1723              :in std_logic_vector(8 DOWNTO 0);
     Lc1724              :in std_logic_vector(8 DOWNTO 0);
     Lc1725              :in std_logic_vector(8 DOWNTO 0);
     Lc1726              :in std_logic_vector(8 DOWNTO 0);
     Lc1727              :in std_logic_vector(8 DOWNTO 0);
     Lc1728              :in std_logic_vector(8 DOWNTO 0);
     Lc1729              :in std_logic_vector(8 DOWNTO 0);
     Lc1730              :in std_logic_vector(8 DOWNTO 0);
     Lc1731              :in std_logic_vector(8 DOWNTO 0);
     Lc1732              :in std_logic_vector(8 DOWNTO 0);
     Lc1733              :in std_logic_vector(8 DOWNTO 0);
     Lc1734              :in std_logic_vector(8 DOWNTO 0);
     Lc1735              :in std_logic_vector(8 DOWNTO 0);
     Lc1736              :in std_logic_vector(8 DOWNTO 0);
     Lc1737              :in std_logic_vector(8 DOWNTO 0);
     Lc1738              :in std_logic_vector(8 DOWNTO 0);
     Lc1739              :in std_logic_vector(8 DOWNTO 0);
     Lc1740              :in std_logic_vector(8 DOWNTO 0);
     Lc1741              :in std_logic_vector(8 DOWNTO 0);
     Lc1742              :in std_logic_vector(8 DOWNTO 0);
     Lc1743              :in std_logic_vector(8 DOWNTO 0);
     Lc1744              :in std_logic_vector(8 DOWNTO 0);
     Lc1745              :in std_logic_vector(8 DOWNTO 0);
     Lc1746              :in std_logic_vector(8 DOWNTO 0);
     Lc1747              :in std_logic_vector(8 DOWNTO 0);
     Lc1748              :in std_logic_vector(8 DOWNTO 0);
     Lc1749              :in std_logic_vector(8 DOWNTO 0);
     Lc1750              :in std_logic_vector(8 DOWNTO 0);
     Lc1751              :in std_logic_vector(8 DOWNTO 0);
     Lc1752              :in std_logic_vector(8 DOWNTO 0);
     Lc1753              :in std_logic_vector(8 DOWNTO 0);
     Lc1754              :in std_logic_vector(8 DOWNTO 0);
     Lc1755              :in std_logic_vector(8 DOWNTO 0);
     Lc1756              :in std_logic_vector(8 DOWNTO 0);
     Lc1757              :in std_logic_vector(8 DOWNTO 0);
     Lc1758              :in std_logic_vector(8 DOWNTO 0);
     Lc1759              :in std_logic_vector(8 DOWNTO 0);
     Lc1760              :in std_logic_vector(8 DOWNTO 0);
     Lc1761              :in std_logic_vector(8 DOWNTO 0);
     Lc1762              :in std_logic_vector(8 DOWNTO 0);
     Lc1763              :in std_logic_vector(8 DOWNTO 0);
     Lc1764              :in std_logic_vector(8 DOWNTO 0);
     Lc1765              :in std_logic_vector(8 DOWNTO 0);
     Lc1766              :in std_logic_vector(8 DOWNTO 0);
     Lc1767              :in std_logic_vector(8 DOWNTO 0);
     Lc1768              :in std_logic_vector(8 DOWNTO 0);
     Lc1769              :in std_logic_vector(8 DOWNTO 0);
     Lc1770              :in std_logic_vector(8 DOWNTO 0);
     Lc1771              :in std_logic_vector(8 DOWNTO 0);
     Lc1772              :in std_logic_vector(8 DOWNTO 0);
     Lc1773              :in std_logic_vector(8 DOWNTO 0);
     Lc1774              :in std_logic_vector(8 DOWNTO 0);
     Lc1775              :in std_logic_vector(8 DOWNTO 0);
     Lc1776              :in std_logic_vector(8 DOWNTO 0);
     Lc1777              :in std_logic_vector(8 DOWNTO 0);
     Lc1778              :in std_logic_vector(8 DOWNTO 0);
     Lc1779              :in std_logic_vector(8 DOWNTO 0);
     Lc1780              :in std_logic_vector(8 DOWNTO 0);
     Lc1781              :in std_logic_vector(8 DOWNTO 0);
     Lc1782              :in std_logic_vector(8 DOWNTO 0);
     Lc1783              :in std_logic_vector(8 DOWNTO 0);
     Lc1784              :in std_logic_vector(8 DOWNTO 0);
     Lc1785              :in std_logic_vector(8 DOWNTO 0);
     Lc1786              :in std_logic_vector(8 DOWNTO 0);
     Lc1787              :in std_logic_vector(8 DOWNTO 0);
     Lc1788              :in std_logic_vector(8 DOWNTO 0);
     Lc1789              :in std_logic_vector(8 DOWNTO 0);
     Lc1790              :in std_logic_vector(8 DOWNTO 0);
     Lc1791              :in std_logic_vector(8 DOWNTO 0);
     Lc1792              :in std_logic_vector(8 DOWNTO 0);
     Lc1793              :in std_logic_vector(8 DOWNTO 0);
     Lc1794              :in std_logic_vector(8 DOWNTO 0);
     Lc1795              :in std_logic_vector(8 DOWNTO 0);
     Lc1796              :in std_logic_vector(8 DOWNTO 0);
     Lc1797              :in std_logic_vector(8 DOWNTO 0);
     Lc1798              :in std_logic_vector(8 DOWNTO 0);
     Lc1799              :in std_logic_vector(8 DOWNTO 0);
     Lc1800              :in std_logic_vector(8 DOWNTO 0);
     Lc1801              :in std_logic_vector(8 DOWNTO 0);
     Lc1802              :in std_logic_vector(8 DOWNTO 0);
     Lc1803              :in std_logic_vector(8 DOWNTO 0);
     Lc1804              :in std_logic_vector(8 DOWNTO 0);
     Lc1805              :in std_logic_vector(8 DOWNTO 0);
     Lc1806              :in std_logic_vector(8 DOWNTO 0);
     Lc1807              :in std_logic_vector(8 DOWNTO 0);
     Lc1808              :in std_logic_vector(8 DOWNTO 0);
     Lc1809              :in std_logic_vector(8 DOWNTO 0);
     Lc1810              :in std_logic_vector(8 DOWNTO 0);
     Lc1811              :in std_logic_vector(8 DOWNTO 0);
     Lc1812              :in std_logic_vector(8 DOWNTO 0);
     Lc1813              :in std_logic_vector(8 DOWNTO 0);
     Lc1814              :in std_logic_vector(8 DOWNTO 0);
     Lc1815              :in std_logic_vector(8 DOWNTO 0);
     Lc1816              :in std_logic_vector(8 DOWNTO 0);
     Lc1817              :in std_logic_vector(8 DOWNTO 0);
     Lc1818              :in std_logic_vector(8 DOWNTO 0);
     Lc1819              :in std_logic_vector(8 DOWNTO 0);
     Lc1820              :in std_logic_vector(8 DOWNTO 0);
     Lc1821              :in std_logic_vector(8 DOWNTO 0);
     Lc1822              :in std_logic_vector(8 DOWNTO 0);
     Lc1823              :in std_logic_vector(8 DOWNTO 0);
     Lc1824              :in std_logic_vector(8 DOWNTO 0);
     Lc1825              :in std_logic_vector(8 DOWNTO 0);
     Lc1826              :in std_logic_vector(8 DOWNTO 0);
     Lc1827              :in std_logic_vector(8 DOWNTO 0);
     Lc1828              :in std_logic_vector(8 DOWNTO 0);
     Lc1829              :in std_logic_vector(8 DOWNTO 0);
     Lc1830              :in std_logic_vector(8 DOWNTO 0);
     Lc1831              :in std_logic_vector(8 DOWNTO 0);
     Lc1832              :in std_logic_vector(8 DOWNTO 0);
     Lc1833              :in std_logic_vector(8 DOWNTO 0);
     Lc1834              :in std_logic_vector(8 DOWNTO 0);
     Lc1835              :in std_logic_vector(8 DOWNTO 0);
     Lc1836              :in std_logic_vector(8 DOWNTO 0);
     Lc1837              :in std_logic_vector(8 DOWNTO 0);
     Lc1838              :in std_logic_vector(8 DOWNTO 0);
     Lc1839              :in std_logic_vector(8 DOWNTO 0);
     Lc1840              :in std_logic_vector(8 DOWNTO 0);
     Lc1841              :in std_logic_vector(8 DOWNTO 0);
     Lc1842              :in std_logic_vector(8 DOWNTO 0);
     Lc1843              :in std_logic_vector(8 DOWNTO 0);
     Lc1844              :in std_logic_vector(8 DOWNTO 0);
     Lc1845              :in std_logic_vector(8 DOWNTO 0);
     Lc1846              :in std_logic_vector(8 DOWNTO 0);
     Lc1847              :in std_logic_vector(8 DOWNTO 0);
     Lc1848              :in std_logic_vector(8 DOWNTO 0);
     Lc1849              :in std_logic_vector(8 DOWNTO 0);
     Lc1850              :in std_logic_vector(8 DOWNTO 0);
     Lc1851              :in std_logic_vector(8 DOWNTO 0);
     Lc1852              :in std_logic_vector(8 DOWNTO 0);
     Lc1853              :in std_logic_vector(8 DOWNTO 0);
     Lc1854              :in std_logic_vector(8 DOWNTO 0);
     Lc1855              :in std_logic_vector(8 DOWNTO 0);
     Lc1856              :in std_logic_vector(8 DOWNTO 0);
     Lc1857              :in std_logic_vector(8 DOWNTO 0);
     Lc1858              :in std_logic_vector(8 DOWNTO 0);
     Lc1859              :in std_logic_vector(8 DOWNTO 0);
     Lc1860              :in std_logic_vector(8 DOWNTO 0);
     Lc1861              :in std_logic_vector(8 DOWNTO 0);
     Lc1862              :in std_logic_vector(8 DOWNTO 0);
     Lc1863              :in std_logic_vector(8 DOWNTO 0);
     Lc1864              :in std_logic_vector(8 DOWNTO 0);
     Lc1865              :in std_logic_vector(8 DOWNTO 0);
     Lc1866              :in std_logic_vector(8 DOWNTO 0);
     Lc1867              :in std_logic_vector(8 DOWNTO 0);
     Lc1868              :in std_logic_vector(8 DOWNTO 0);
     Lc1869              :in std_logic_vector(8 DOWNTO 0);
     Lc1870              :in std_logic_vector(8 DOWNTO 0);
     Lc1871              :in std_logic_vector(8 DOWNTO 0);
     Lc1872              :in std_logic_vector(8 DOWNTO 0);
     Lc1873              :in std_logic_vector(8 DOWNTO 0);
     Lc1874              :in std_logic_vector(8 DOWNTO 0);
     Lc1875              :in std_logic_vector(8 DOWNTO 0);
     Lc1876              :in std_logic_vector(8 DOWNTO 0);
     Lc1877              :in std_logic_vector(8 DOWNTO 0);
     Lc1878              :in std_logic_vector(8 DOWNTO 0);
     Lc1879              :in std_logic_vector(8 DOWNTO 0);
     Lc1880              :in std_logic_vector(8 DOWNTO 0);
     Lc1881              :in std_logic_vector(8 DOWNTO 0);
     Lc1882              :in std_logic_vector(8 DOWNTO 0);
     Lc1883              :in std_logic_vector(8 DOWNTO 0);
     Lc1884              :in std_logic_vector(8 DOWNTO 0);
     Lc1885              :in std_logic_vector(8 DOWNTO 0);
     Lc1886              :in std_logic_vector(8 DOWNTO 0);
     Lc1887              :in std_logic_vector(8 DOWNTO 0);
     Lc1888              :in std_logic_vector(8 DOWNTO 0);
     Lc1889              :in std_logic_vector(8 DOWNTO 0);
     Lc1890              :in std_logic_vector(8 DOWNTO 0);
     Lc1891              :in std_logic_vector(8 DOWNTO 0);
     Lc1892              :in std_logic_vector(8 DOWNTO 0);
     Lc1893              :in std_logic_vector(8 DOWNTO 0);
     Lc1894              :in std_logic_vector(8 DOWNTO 0);
     Lc1895              :in std_logic_vector(8 DOWNTO 0);
     Lc1896              :in std_logic_vector(8 DOWNTO 0);
     Lc1897              :in std_logic_vector(8 DOWNTO 0);
     Lc1898              :in std_logic_vector(8 DOWNTO 0);
     Lc1899              :in std_logic_vector(8 DOWNTO 0);
     Lc1900              :in std_logic_vector(8 DOWNTO 0);
     Lc1901              :in std_logic_vector(8 DOWNTO 0);
     Lc1902              :in std_logic_vector(8 DOWNTO 0);
     Lc1903              :in std_logic_vector(8 DOWNTO 0);
     Lc1904              :in std_logic_vector(8 DOWNTO 0);
     Lc1905              :in std_logic_vector(8 DOWNTO 0);
     Lc1906              :in std_logic_vector(8 DOWNTO 0);
     Lc1907              :in std_logic_vector(8 DOWNTO 0);
     Lc1908              :in std_logic_vector(8 DOWNTO 0);
     Lc1909              :in std_logic_vector(8 DOWNTO 0);
     Lc1910              :in std_logic_vector(8 DOWNTO 0);
     Lc1911              :in std_logic_vector(8 DOWNTO 0);
     Lc1912              :in std_logic_vector(8 DOWNTO 0);
     Lc1913              :in std_logic_vector(8 DOWNTO 0);
     Lc1914              :in std_logic_vector(8 DOWNTO 0);
     Lc1915              :in std_logic_vector(8 DOWNTO 0);
     Lc1916              :in std_logic_vector(8 DOWNTO 0);
     Lc1917              :in std_logic_vector(8 DOWNTO 0);
     Lc1918              :in std_logic_vector(8 DOWNTO 0);
     Lc1919              :in std_logic_vector(8 DOWNTO 0);
     Lc1920              :in std_logic_vector(8 DOWNTO 0);
     Lc1921              :in std_logic_vector(8 DOWNTO 0);
     Lc1922              :in std_logic_vector(8 DOWNTO 0);
     Lc1923              :in std_logic_vector(8 DOWNTO 0);
     Lc1924              :in std_logic_vector(8 DOWNTO 0);
     Lc1925              :in std_logic_vector(8 DOWNTO 0);
     Lc1926              :in std_logic_vector(8 DOWNTO 0);
     Lc1927              :in std_logic_vector(8 DOWNTO 0);
     Lc1928              :in std_logic_vector(8 DOWNTO 0);
     Lc1929              :in std_logic_vector(8 DOWNTO 0);
     Lc1930              :in std_logic_vector(8 DOWNTO 0);
     Lc1931              :in std_logic_vector(8 DOWNTO 0);
     Lc1932              :in std_logic_vector(8 DOWNTO 0);
     Lc1933              :in std_logic_vector(8 DOWNTO 0);
     Lc1934              :in std_logic_vector(8 DOWNTO 0);
     Lc1935              :in std_logic_vector(8 DOWNTO 0);
     Lc1936              :in std_logic_vector(8 DOWNTO 0);
     Lc1937              :in std_logic_vector(8 DOWNTO 0);
     Lc1938              :in std_logic_vector(8 DOWNTO 0);
     Lc1939              :in std_logic_vector(8 DOWNTO 0);
     Lc1940              :in std_logic_vector(8 DOWNTO 0);
     Lc1941              :in std_logic_vector(8 DOWNTO 0);
     Lc1942              :in std_logic_vector(8 DOWNTO 0);
     Lc1943              :in std_logic_vector(8 DOWNTO 0);
     Lc1944              :in std_logic_vector(8 DOWNTO 0);
     Lc1945              :in std_logic_vector(8 DOWNTO 0);
     Lc1946              :in std_logic_vector(8 DOWNTO 0);
     Lc1947              :in std_logic_vector(8 DOWNTO 0);
     Lc1948              :in std_logic_vector(8 DOWNTO 0);
     Lc1949              :in std_logic_vector(8 DOWNTO 0);
     Lc1950              :in std_logic_vector(8 DOWNTO 0);
     Lc1951              :in std_logic_vector(8 DOWNTO 0);
     Lc1952              :in std_logic_vector(8 DOWNTO 0);
     Lc1953              :in std_logic_vector(8 DOWNTO 0);
     Lc1954              :in std_logic_vector(8 DOWNTO 0);
     Lc1955              :in std_logic_vector(8 DOWNTO 0);
     Lc1956              :in std_logic_vector(8 DOWNTO 0);
     Lc1957              :in std_logic_vector(8 DOWNTO 0);
     Lc1958              :in std_logic_vector(8 DOWNTO 0);
     Lc1959              :in std_logic_vector(8 DOWNTO 0);
     Lc1960              :in std_logic_vector(8 DOWNTO 0);
     Lc1961              :in std_logic_vector(8 DOWNTO 0);
     Lc1962              :in std_logic_vector(8 DOWNTO 0);
     Lc1963              :in std_logic_vector(8 DOWNTO 0);
     Lc1964              :in std_logic_vector(8 DOWNTO 0);
     Lc1965              :in std_logic_vector(8 DOWNTO 0);
     Lc1966              :in std_logic_vector(8 DOWNTO 0);
     Lc1967              :in std_logic_vector(8 DOWNTO 0);
     Lc1968              :in std_logic_vector(8 DOWNTO 0);
     Lc1969              :in std_logic_vector(8 DOWNTO 0);
     Lc1970              :in std_logic_vector(8 DOWNTO 0);
     Lc1971              :in std_logic_vector(8 DOWNTO 0);
     Lc1972              :in std_logic_vector(8 DOWNTO 0);
     Lc1973              :in std_logic_vector(8 DOWNTO 0);
     Lc1974              :in std_logic_vector(8 DOWNTO 0);
     Lc1975              :in std_logic_vector(8 DOWNTO 0);
     Lc1976              :in std_logic_vector(8 DOWNTO 0);
     Lc1977              :in std_logic_vector(8 DOWNTO 0);
     Lc1978              :in std_logic_vector(8 DOWNTO 0);
     Lc1979              :in std_logic_vector(8 DOWNTO 0);
     Lc1980              :in std_logic_vector(8 DOWNTO 0);
     Lc1981              :in std_logic_vector(8 DOWNTO 0);
     Lc1982              :in std_logic_vector(8 DOWNTO 0);
     Lc1983              :in std_logic_vector(8 DOWNTO 0);
     Lc1984              :in std_logic_vector(8 DOWNTO 0);
     Lc1985              :in std_logic_vector(8 DOWNTO 0);
     Lc1986              :in std_logic_vector(8 DOWNTO 0);
     Lc1987              :in std_logic_vector(8 DOWNTO 0);
     Lc1988              :in std_logic_vector(8 DOWNTO 0);
     Lc1989              :in std_logic_vector(8 DOWNTO 0);
     Lc1990              :in std_logic_vector(8 DOWNTO 0);
     Lc1991              :in std_logic_vector(8 DOWNTO 0);
     Lc1992              :in std_logic_vector(8 DOWNTO 0);
     Lc1993              :in std_logic_vector(8 DOWNTO 0);
     Lc1994              :in std_logic_vector(8 DOWNTO 0);
     Lc1995              :in std_logic_vector(8 DOWNTO 0);
     Lc1996              :in std_logic_vector(8 DOWNTO 0);
     Lc1997              :in std_logic_vector(8 DOWNTO 0);
     Lc1998              :in std_logic_vector(8 DOWNTO 0);
     Lc1999              :in std_logic_vector(8 DOWNTO 0);
     Lc2000              :in std_logic_vector(8 DOWNTO 0);
     Lc2001              :in std_logic_vector(8 DOWNTO 0);
     Lc2002              :in std_logic_vector(8 DOWNTO 0);
     Lc2003              :in std_logic_vector(8 DOWNTO 0);
     Lc2004              :in std_logic_vector(8 DOWNTO 0);
     Lc2005              :in std_logic_vector(8 DOWNTO 0);
     Lc2006              :in std_logic_vector(8 DOWNTO 0);
     Lc2007              :in std_logic_vector(8 DOWNTO 0);
     Lc2008              :in std_logic_vector(8 DOWNTO 0);
     Lc2009              :in std_logic_vector(8 DOWNTO 0);
     Lc2010              :in std_logic_vector(8 DOWNTO 0);
     Lc2011              :in std_logic_vector(8 DOWNTO 0);
     Lc2012              :in std_logic_vector(8 DOWNTO 0);
     Lc2013              :in std_logic_vector(8 DOWNTO 0);
     Lc2014              :in std_logic_vector(8 DOWNTO 0);
     Lc2015              :in std_logic_vector(8 DOWNTO 0);
     Lc2016              :in std_logic_vector(8 DOWNTO 0);
     Lc2017              :in std_logic_vector(8 DOWNTO 0);
     Lc2018              :in std_logic_vector(8 DOWNTO 0);
     Lc2019              :in std_logic_vector(8 DOWNTO 0);
     Lc2020              :in std_logic_vector(8 DOWNTO 0);
     Lc2021              :in std_logic_vector(8 DOWNTO 0);
     Lc2022              :in std_logic_vector(8 DOWNTO 0);
     Lc2023              :in std_logic_vector(8 DOWNTO 0);
     Lc2024              :in std_logic_vector(8 DOWNTO 0);
     Lc2025              :in std_logic_vector(8 DOWNTO 0);
     Lc2026              :in std_logic_vector(8 DOWNTO 0);
     Lc2027              :in std_logic_vector(8 DOWNTO 0);
     Lc2028              :in std_logic_vector(8 DOWNTO 0);
     Lc2029              :in std_logic_vector(8 DOWNTO 0);
     Lc2030              :in std_logic_vector(8 DOWNTO 0);
     Lc2031              :in std_logic_vector(8 DOWNTO 0);
     Lc2032              :in std_logic_vector(8 DOWNTO 0);
     Lc2033              :in std_logic_vector(8 DOWNTO 0);
     Lc2034              :in std_logic_vector(8 DOWNTO 0);
     Lc2035              :in std_logic_vector(8 DOWNTO 0);
     Lc2036              :in std_logic_vector(8 DOWNTO 0);
     Lc2037              :in std_logic_vector(8 DOWNTO 0);
     Lc2038              :in std_logic_vector(8 DOWNTO 0);
     Lc2039              :in std_logic_vector(8 DOWNTO 0);
     Lc2040              :in std_logic_vector(8 DOWNTO 0);
     Lc2041              :in std_logic_vector(8 DOWNTO 0);
     Lc2042              :in std_logic_vector(8 DOWNTO 0);
     Lc2043              :in std_logic_vector(8 DOWNTO 0);
     Lc2044              :in std_logic_vector(8 DOWNTO 0);
     Lc2045              :in std_logic_vector(8 DOWNTO 0);
     Lc2046              :in std_logic_vector(8 DOWNTO 0);
     Lc2047              :in std_logic_vector(8 DOWNTO 0);
     Lc2048              :in std_logic_vector(8 DOWNTO 0);
     Lc2049              :in std_logic_vector(8 DOWNTO 0);
     Lc2050              :in std_logic_vector(8 DOWNTO 0);
     Lc2051              :in std_logic_vector(8 DOWNTO 0);
     Lc2052              :in std_logic_vector(8 DOWNTO 0);
     Lc2053              :in std_logic_vector(8 DOWNTO 0);
     Lc2054              :in std_logic_vector(8 DOWNTO 0);
     Lc2055              :in std_logic_vector(8 DOWNTO 0);
     Lc2056              :in std_logic_vector(8 DOWNTO 0);
     Lc2057              :in std_logic_vector(8 DOWNTO 0);
     Lc2058              :in std_logic_vector(8 DOWNTO 0);
     Lc2059              :in std_logic_vector(8 DOWNTO 0);
     Lc2060              :in std_logic_vector(8 DOWNTO 0);
     Lc2061              :in std_logic_vector(8 DOWNTO 0);
     Lc2062              :in std_logic_vector(8 DOWNTO 0);
     Lc2063              :in std_logic_vector(8 DOWNTO 0);
     Lc2064              :in std_logic_vector(8 DOWNTO 0);
     Lc2065              :in std_logic_vector(8 DOWNTO 0);
     Lc2066              :in std_logic_vector(8 DOWNTO 0);
     Lc2067              :in std_logic_vector(8 DOWNTO 0);
     Lc2068              :in std_logic_vector(8 DOWNTO 0);
     Lc2069              :in std_logic_vector(8 DOWNTO 0);
     Lc2070              :in std_logic_vector(8 DOWNTO 0);
     Lc2071              :in std_logic_vector(8 DOWNTO 0);
     Lc2072              :in std_logic_vector(8 DOWNTO 0);
     Lc2073              :in std_logic_vector(8 DOWNTO 0);
     Lc2074              :in std_logic_vector(8 DOWNTO 0);
     Lc2075              :in std_logic_vector(8 DOWNTO 0);
     Lc2076              :in std_logic_vector(8 DOWNTO 0);
     Lc2077              :in std_logic_vector(8 DOWNTO 0);
     Lc2078              :in std_logic_vector(8 DOWNTO 0);
     Lc2079              :in std_logic_vector(8 DOWNTO 0);
     Lc2080              :in std_logic_vector(8 DOWNTO 0);
     Lc2081              :in std_logic_vector(8 DOWNTO 0);
     Lc2082              :in std_logic_vector(8 DOWNTO 0);
     Lc2083              :in std_logic_vector(8 DOWNTO 0);
     Lc2084              :in std_logic_vector(8 DOWNTO 0);
     Lc2085              :in std_logic_vector(8 DOWNTO 0);
     Lc2086              :in std_logic_vector(8 DOWNTO 0);
     Lc2087              :in std_logic_vector(8 DOWNTO 0);
     Lc2088              :in std_logic_vector(8 DOWNTO 0);
     Lc2089              :in std_logic_vector(8 DOWNTO 0);
     Lc2090              :in std_logic_vector(8 DOWNTO 0);
     Lc2091              :in std_logic_vector(8 DOWNTO 0);
     Lc2092              :in std_logic_vector(8 DOWNTO 0);
     Lc2093              :in std_logic_vector(8 DOWNTO 0);
     Lc2094              :in std_logic_vector(8 DOWNTO 0);
     Lc2095              :in std_logic_vector(8 DOWNTO 0);
     Lc2096              :in std_logic_vector(8 DOWNTO 0);
     Lc2097              :in std_logic_vector(8 DOWNTO 0);
     Lc2098              :in std_logic_vector(8 DOWNTO 0);
     Lc2099              :in std_logic_vector(8 DOWNTO 0);
     Lc2100              :in std_logic_vector(8 DOWNTO 0);
     Lc2101              :in std_logic_vector(8 DOWNTO 0);
     Lc2102              :in std_logic_vector(8 DOWNTO 0);
     Lc2103              :in std_logic_vector(8 DOWNTO 0);
     Lc2104              :in std_logic_vector(8 DOWNTO 0);
     Lc2105              :in std_logic_vector(8 DOWNTO 0);
     Lc2106              :in std_logic_vector(8 DOWNTO 0);
     Lc2107              :in std_logic_vector(8 DOWNTO 0);
     Lc2108              :in std_logic_vector(8 DOWNTO 0);
     Lc2109              :in std_logic_vector(8 DOWNTO 0);
     Lc2110              :in std_logic_vector(8 DOWNTO 0);
     Lc2111              :in std_logic_vector(8 DOWNTO 0);
     Lc2112              :in std_logic_vector(8 DOWNTO 0);
     Lc2113              :in std_logic_vector(8 DOWNTO 0);
     Lc2114              :in std_logic_vector(8 DOWNTO 0);
     Lc2115              :in std_logic_vector(8 DOWNTO 0);
     Lc2116              :in std_logic_vector(8 DOWNTO 0);
     Lc2117              :in std_logic_vector(8 DOWNTO 0);
     Lc2118              :in std_logic_vector(8 DOWNTO 0);
     Lc2119              :in std_logic_vector(8 DOWNTO 0);
     Lc2120              :in std_logic_vector(8 DOWNTO 0);
     Lc2121              :in std_logic_vector(8 DOWNTO 0);
     Lc2122              :in std_logic_vector(8 DOWNTO 0);
     Lc2123              :in std_logic_vector(8 DOWNTO 0);
     Lc2124              :in std_logic_vector(8 DOWNTO 0);
     Lc2125              :in std_logic_vector(8 DOWNTO 0);
     Lc2126              :in std_logic_vector(8 DOWNTO 0);
     Lc2127              :in std_logic_vector(8 DOWNTO 0);
     Lc2128              :in std_logic_vector(8 DOWNTO 0);
     Lc2129              :in std_logic_vector(8 DOWNTO 0);
     Lc2130              :in std_logic_vector(8 DOWNTO 0);
     Lc2131              :in std_logic_vector(8 DOWNTO 0);
     Lc2132              :in std_logic_vector(8 DOWNTO 0);
     Lc2133              :in std_logic_vector(8 DOWNTO 0);
     Lc2134              :in std_logic_vector(8 DOWNTO 0);
     Lc2135              :in std_logic_vector(8 DOWNTO 0);
     Lc2136              :in std_logic_vector(8 DOWNTO 0);
     Lc2137              :in std_logic_vector(8 DOWNTO 0);
     Lc2138              :in std_logic_vector(8 DOWNTO 0);
     Lc2139              :in std_logic_vector(8 DOWNTO 0);
     Lc2140              :in std_logic_vector(8 DOWNTO 0);
     Lc2141              :in std_logic_vector(8 DOWNTO 0);
     Lc2142              :in std_logic_vector(8 DOWNTO 0);
     Lc2143              :in std_logic_vector(8 DOWNTO 0);
     Lc2144              :in std_logic_vector(8 DOWNTO 0);
     Lc2145              :in std_logic_vector(8 DOWNTO 0);
     Lc2146              :in std_logic_vector(8 DOWNTO 0);
     Lc2147              :in std_logic_vector(8 DOWNTO 0);
     Lc2148              :in std_logic_vector(8 DOWNTO 0);
     Lc2149              :in std_logic_vector(8 DOWNTO 0);
     Lc2150              :in std_logic_vector(8 DOWNTO 0);
     Lc2151              :in std_logic_vector(8 DOWNTO 0);
     Lc2152              :in std_logic_vector(8 DOWNTO 0);
     Lc2153              :in std_logic_vector(8 DOWNTO 0);
     Lc2154              :in std_logic_vector(8 DOWNTO 0);
     Lc2155              :in std_logic_vector(8 DOWNTO 0);
     Lc2156              :in std_logic_vector(8 DOWNTO 0);
     Lc2157              :in std_logic_vector(8 DOWNTO 0);
     Lc2158              :in std_logic_vector(8 DOWNTO 0);
     Lc2159              :in std_logic_vector(8 DOWNTO 0);
     Lc2160              :in std_logic_vector(8 DOWNTO 0);
     Lc2161              :in std_logic_vector(8 DOWNTO 0);
     Lc2162              :in std_logic_vector(8 DOWNTO 0);
     Lc2163              :in std_logic_vector(8 DOWNTO 0);
     Lc2164              :in std_logic_vector(8 DOWNTO 0);
     Lc2165              :in std_logic_vector(8 DOWNTO 0);
     Lc2166              :in std_logic_vector(8 DOWNTO 0);
     Lc2167              :in std_logic_vector(8 DOWNTO 0);
     Lc2168              :in std_logic_vector(8 DOWNTO 0);
     Lc2169              :in std_logic_vector(8 DOWNTO 0);
     Lc2170              :in std_logic_vector(8 DOWNTO 0);
     Lc2171              :in std_logic_vector(8 DOWNTO 0);
     Lc2172              :in std_logic_vector(8 DOWNTO 0);
     Lc2173              :in std_logic_vector(8 DOWNTO 0);
     Lc2174              :in std_logic_vector(8 DOWNTO 0);
     Lc2175              :in std_logic_vector(8 DOWNTO 0);
     Lc2176              :in std_logic_vector(8 DOWNTO 0);
     Lc2177              :in std_logic_vector(8 DOWNTO 0);
     Lc2178              :in std_logic_vector(8 DOWNTO 0);
     Lc2179              :in std_logic_vector(8 DOWNTO 0);
     Lc2180              :in std_logic_vector(8 DOWNTO 0);
     Lc2181              :in std_logic_vector(8 DOWNTO 0);
     Lc2182              :in std_logic_vector(8 DOWNTO 0);
     Lc2183              :in std_logic_vector(8 DOWNTO 0);
     Lc2184              :in std_logic_vector(8 DOWNTO 0);
     Lc2185              :in std_logic_vector(8 DOWNTO 0);
     Lc2186              :in std_logic_vector(8 DOWNTO 0);
     Lc2187              :in std_logic_vector(8 DOWNTO 0);
     Lc2188              :in std_logic_vector(8 DOWNTO 0);
     Lc2189              :in std_logic_vector(8 DOWNTO 0);
     Lc2190              :in std_logic_vector(8 DOWNTO 0);
     Lc2191              :in std_logic_vector(8 DOWNTO 0);
     Lc2192              :in std_logic_vector(8 DOWNTO 0);
     Lc2193              :in std_logic_vector(8 DOWNTO 0);
     Lc2194              :in std_logic_vector(8 DOWNTO 0);
     Lc2195              :in std_logic_vector(8 DOWNTO 0);
     Lc2196              :in std_logic_vector(8 DOWNTO 0);
     Lc2197              :in std_logic_vector(8 DOWNTO 0);
     Lc2198              :in std_logic_vector(8 DOWNTO 0);
     Lc2199              :in std_logic_vector(8 DOWNTO 0);
     Lc2200              :in std_logic_vector(8 DOWNTO 0);
     Lc2201              :in std_logic_vector(8 DOWNTO 0);
     Lc2202              :in std_logic_vector(8 DOWNTO 0);
     Lc2203              :in std_logic_vector(8 DOWNTO 0);
     Lc2204              :in std_logic_vector(8 DOWNTO 0);
     Lc2205              :in std_logic_vector(8 DOWNTO 0);
     Lc2206              :in std_logic_vector(8 DOWNTO 0);
     Lc2207              :in std_logic_vector(8 DOWNTO 0);
     Lc2208              :in std_logic_vector(8 DOWNTO 0);
     Lc2209              :in std_logic_vector(8 DOWNTO 0);
     Lc2210              :in std_logic_vector(8 DOWNTO 0);
     Lc2211              :in std_logic_vector(8 DOWNTO 0);
     Lc2212              :in std_logic_vector(8 DOWNTO 0);
     Lc2213              :in std_logic_vector(8 DOWNTO 0);
     Lc2214              :in std_logic_vector(8 DOWNTO 0);
     Lc2215              :in std_logic_vector(8 DOWNTO 0);
     Lc2216              :in std_logic_vector(8 DOWNTO 0);
     Lc2217              :in std_logic_vector(8 DOWNTO 0);
     Lc2218              :in std_logic_vector(8 DOWNTO 0);
     Lc2219              :in std_logic_vector(8 DOWNTO 0);
     Lc2220              :in std_logic_vector(8 DOWNTO 0);
     Lc2221              :in std_logic_vector(8 DOWNTO 0);
     Lc2222              :in std_logic_vector(8 DOWNTO 0);
     Lc2223              :in std_logic_vector(8 DOWNTO 0);
     Lc2224              :in std_logic_vector(8 DOWNTO 0);
     Lc2225              :in std_logic_vector(8 DOWNTO 0);
     Lc2226              :in std_logic_vector(8 DOWNTO 0);
     Lc2227              :in std_logic_vector(8 DOWNTO 0);
     Lc2228              :in std_logic_vector(8 DOWNTO 0);
     Lc2229              :in std_logic_vector(8 DOWNTO 0);
     Lc2230              :in std_logic_vector(8 DOWNTO 0);
     Lc2231              :in std_logic_vector(8 DOWNTO 0);
     Lc2232              :in std_logic_vector(8 DOWNTO 0);
     Lc2233              :in std_logic_vector(8 DOWNTO 0);
     Lc2234              :in std_logic_vector(8 DOWNTO 0);
     Lc2235              :in std_logic_vector(8 DOWNTO 0);
     Lc2236              :in std_logic_vector(8 DOWNTO 0);
     Lc2237              :in std_logic_vector(8 DOWNTO 0);
     Lc2238              :in std_logic_vector(8 DOWNTO 0);
     Lc2239              :in std_logic_vector(8 DOWNTO 0);
     Lc2240              :in std_logic_vector(8 DOWNTO 0);
     Lc2241              :in std_logic_vector(8 DOWNTO 0);
     Lc2242              :in std_logic_vector(8 DOWNTO 0);
     Lc2243              :in std_logic_vector(8 DOWNTO 0);
     Lc2244              :in std_logic_vector(8 DOWNTO 0);
     Lc2245              :in std_logic_vector(8 DOWNTO 0);
     Lc2246              :in std_logic_vector(8 DOWNTO 0);
     Lc2247              :in std_logic_vector(8 DOWNTO 0);
     Lc2248              :in std_logic_vector(8 DOWNTO 0);
     Lc2249              :in std_logic_vector(8 DOWNTO 0);
     Lc2250              :in std_logic_vector(8 DOWNTO 0);
     Lc2251              :in std_logic_vector(8 DOWNTO 0);
     Lc2252              :in std_logic_vector(8 DOWNTO 0);
     Lc2253              :in std_logic_vector(8 DOWNTO 0);
     Lc2254              :in std_logic_vector(8 DOWNTO 0);
     Lc2255              :in std_logic_vector(8 DOWNTO 0);
     Lc2256              :in std_logic_vector(8 DOWNTO 0);
     Lc2257              :in std_logic_vector(8 DOWNTO 0);
     Lc2258              :in std_logic_vector(8 DOWNTO 0);
     Lc2259              :in std_logic_vector(8 DOWNTO 0);
     Lc2260              :in std_logic_vector(8 DOWNTO 0);
     Lc2261              :in std_logic_vector(8 DOWNTO 0);
     Lc2262              :in std_logic_vector(8 DOWNTO 0);
     Lc2263              :in std_logic_vector(8 DOWNTO 0);
     Lc2264              :in std_logic_vector(8 DOWNTO 0);
     Lc2265              :in std_logic_vector(8 DOWNTO 0);
     Lc2266              :in std_logic_vector(8 DOWNTO 0);
     Lc2267              :in std_logic_vector(8 DOWNTO 0);
     Lc2268              :in std_logic_vector(8 DOWNTO 0);
     Lc2269              :in std_logic_vector(8 DOWNTO 0);
     Lc2270              :in std_logic_vector(8 DOWNTO 0);
     Lc2271              :in std_logic_vector(8 DOWNTO 0);
     Lc2272              :in std_logic_vector(8 DOWNTO 0);
     Lc2273              :in std_logic_vector(8 DOWNTO 0);
     Lc2274              :in std_logic_vector(8 DOWNTO 0);
     Lc2275              :in std_logic_vector(8 DOWNTO 0);
     Lc2276              :in std_logic_vector(8 DOWNTO 0);
     Lc2277              :in std_logic_vector(8 DOWNTO 0);
     Lc2278              :in std_logic_vector(8 DOWNTO 0);
     Lc2279              :in std_logic_vector(8 DOWNTO 0);
     Lc2280              :in std_logic_vector(8 DOWNTO 0);
     Lc2281              :in std_logic_vector(8 DOWNTO 0);
     Lc2282              :in std_logic_vector(8 DOWNTO 0);
     Lc2283              :in std_logic_vector(8 DOWNTO 0);
     Lc2284              :in std_logic_vector(8 DOWNTO 0);
     Lc2285              :in std_logic_vector(8 DOWNTO 0);
     Lc2286              :in std_logic_vector(8 DOWNTO 0);
     Lc2287              :in std_logic_vector(8 DOWNTO 0);
     Lc2288              :in std_logic_vector(8 DOWNTO 0);
     Lc2289              :in std_logic_vector(8 DOWNTO 0);
     Lc2290              :in std_logic_vector(8 DOWNTO 0);
     Lc2291              :in std_logic_vector(8 DOWNTO 0);
     Lc2292              :in std_logic_vector(8 DOWNTO 0);
     Lc2293              :in std_logic_vector(8 DOWNTO 0);
     Lc2294              :in std_logic_vector(8 DOWNTO 0);
     Lc2295              :in std_logic_vector(8 DOWNTO 0);
     Lc2296              :in std_logic_vector(8 DOWNTO 0);
     Lc2297              :in std_logic_vector(8 DOWNTO 0);
     Lc2298              :in std_logic_vector(8 DOWNTO 0);
     Lc2299              :in std_logic_vector(8 DOWNTO 0);
     Lc2300              :in std_logic_vector(8 DOWNTO 0);
     Lc2301              :in std_logic_vector(8 DOWNTO 0);
     Lc2302              :in std_logic_vector(8 DOWNTO 0);
     Lc2303              :in std_logic_vector(8 DOWNTO 0);
     Lc2304              :in std_logic_vector(8 DOWNTO 0);
     out1            :out std_logic;
     out2            :out std_logic;
     out3            :out std_logic;
     out4            :out std_logic;
     out5            :out std_logic;
     out6            :out std_logic;
     out7            :out std_logic;
     out8            :out std_logic;
     out9            :out std_logic;
     out10            :out std_logic;
     out11            :out std_logic;
     out12            :out std_logic;
     out13            :out std_logic;
     out14            :out std_logic;
     out15            :out std_logic;
     out16            :out std_logic;
     out17            :out std_logic;
     out18            :out std_logic;
     out19            :out std_logic;
     out20            :out std_logic;
     out21            :out std_logic;
     out22            :out std_logic;
     out23            :out std_logic;
     out24            :out std_logic;
     out25            :out std_logic;
     out26            :out std_logic;
     out27            :out std_logic;
     out28            :out std_logic;
     out29            :out std_logic;
     out30            :out std_logic;
     out31            :out std_logic;
     out32            :out std_logic;
     out33            :out std_logic;
     out34            :out std_logic;
     out35            :out std_logic;
     out36            :out std_logic;
     out37            :out std_logic;
     out38            :out std_logic;
     out39            :out std_logic;
     out40            :out std_logic;
     out41            :out std_logic;
     out42            :out std_logic;
     out43            :out std_logic;
     out44            :out std_logic;
     out45            :out std_logic;
     out46            :out std_logic;
     out47            :out std_logic;
     out48            :out std_logic;
     out49            :out std_logic;
     out50            :out std_logic;
     out51            :out std_logic;
     out52            :out std_logic;
     out53            :out std_logic;
     out54            :out std_logic;
     out55            :out std_logic;
     out56            :out std_logic;
     out57            :out std_logic;
     out58            :out std_logic;
     out59            :out std_logic;
     out60            :out std_logic;
     out61            :out std_logic;
     out62            :out std_logic;
     out63            :out std_logic;
     out64            :out std_logic;
     out65            :out std_logic;
     out66            :out std_logic;
     out67            :out std_logic;
     out68            :out std_logic;
     out69            :out std_logic;
     out70            :out std_logic;
     out71            :out std_logic;
     out72            :out std_logic;
     out73            :out std_logic;
     out74            :out std_logic;
     out75            :out std_logic;
     out76            :out std_logic;
     out77            :out std_logic;
     out78            :out std_logic;
     out79            :out std_logic;
     out80            :out std_logic;
     out81            :out std_logic;
     out82            :out std_logic;
     out83            :out std_logic;
     out84            :out std_logic;
     out85            :out std_logic;
     out86            :out std_logic;
     out87            :out std_logic;
     out88            :out std_logic;
     out89            :out std_logic;
     out90            :out std_logic;
     out91            :out std_logic;
     out92            :out std_logic;
     out93            :out std_logic;
     out94            :out std_logic;
     out95            :out std_logic;
     out96            :out std_logic;
     out97            :out std_logic;
     out98            :out std_logic;
     out99            :out std_logic;
     out100            :out std_logic;
     out101            :out std_logic;
     out102            :out std_logic;
     out103            :out std_logic;
     out104            :out std_logic;
     out105            :out std_logic;
     out106            :out std_logic;
     out107            :out std_logic;
     out108            :out std_logic;
     out109            :out std_logic;
     out110            :out std_logic;
     out111            :out std_logic;
     out112            :out std_logic;
     out113            :out std_logic;
     out114            :out std_logic;
     out115            :out std_logic;
     out116            :out std_logic;
     out117            :out std_logic;
     out118            :out std_logic;
     out119            :out std_logic;
     out120            :out std_logic;
     out121            :out std_logic;
     out122            :out std_logic;
     out123            :out std_logic;
     out124            :out std_logic;
     out125            :out std_logic;
     out126            :out std_logic;
     out127            :out std_logic;
     out128            :out std_logic;
     out129            :out std_logic;
     out130            :out std_logic;
     out131            :out std_logic;
     out132            :out std_logic;
     out133            :out std_logic;
     out134            :out std_logic;
     out135            :out std_logic;
     out136            :out std_logic;
     out137            :out std_logic;
     out138            :out std_logic;
     out139            :out std_logic;
     out140            :out std_logic;
     out141            :out std_logic;
     out142            :out std_logic;
     out143            :out std_logic;
     out144            :out std_logic;
     out145            :out std_logic;
     out146            :out std_logic;
     out147            :out std_logic;
     out148            :out std_logic;
     out149            :out std_logic;
     out150            :out std_logic;
     out151            :out std_logic;
     out152            :out std_logic;
     out153            :out std_logic;
     out154            :out std_logic;
     out155            :out std_logic;
     out156            :out std_logic;
     out157            :out std_logic;
     out158            :out std_logic;
     out159            :out std_logic;
     out160            :out std_logic;
     out161            :out std_logic;
     out162            :out std_logic;
     out163            :out std_logic;
     out164            :out std_logic;
     out165            :out std_logic;
     out166            :out std_logic;
     out167            :out std_logic;
     out168            :out std_logic;
     out169            :out std_logic;
     out170            :out std_logic;
     out171            :out std_logic;
     out172            :out std_logic;
     out173            :out std_logic;
     out174            :out std_logic;
     out175            :out std_logic;
     out176            :out std_logic;
     out177            :out std_logic;
     out178            :out std_logic;
     out179            :out std_logic;
     out180            :out std_logic;
     out181            :out std_logic;
     out182            :out std_logic;
     out183            :out std_logic;
     out184            :out std_logic;
     out185            :out std_logic;
     out186            :out std_logic;
     out187            :out std_logic;
     out188            :out std_logic;
     out189            :out std_logic;
     out190            :out std_logic;
     out191            :out std_logic;
     out192            :out std_logic;
     out193            :out std_logic;
     out194            :out std_logic;
     out195            :out std_logic;
     out196            :out std_logic;
     out197            :out std_logic;
     out198            :out std_logic;
     out199            :out std_logic;
     out200            :out std_logic;
     out201            :out std_logic;
     out202            :out std_logic;
     out203            :out std_logic;
     out204            :out std_logic;
     out205            :out std_logic;
     out206            :out std_logic;
     out207            :out std_logic;
     out208            :out std_logic;
     out209            :out std_logic;
     out210            :out std_logic;
     out211            :out std_logic;
     out212            :out std_logic;
     out213            :out std_logic;
     out214            :out std_logic;
     out215            :out std_logic;
     out216            :out std_logic;
     out217            :out std_logic;
     out218            :out std_logic;
     out219            :out std_logic;
     out220            :out std_logic;
     out221            :out std_logic;
     out222            :out std_logic;
     out223            :out std_logic;
     out224            :out std_logic;
     out225            :out std_logic;
     out226            :out std_logic;
     out227            :out std_logic;
     out228            :out std_logic;
     out229            :out std_logic;
     out230            :out std_logic;
     out231            :out std_logic;
     out232            :out std_logic;
     out233            :out std_logic;
     out234            :out std_logic;
     out235            :out std_logic;
     out236            :out std_logic;
     out237            :out std_logic;
     out238            :out std_logic;
     out239            :out std_logic;
     out240            :out std_logic;
     out241            :out std_logic;
     out242            :out std_logic;
     out243            :out std_logic;
     out244            :out std_logic;
     out245            :out std_logic;
     out246            :out std_logic;
     out247            :out std_logic;
     out248            :out std_logic;
     out249            :out std_logic;
     out250            :out std_logic;
     out251            :out std_logic;
     out252            :out std_logic;
     out253            :out std_logic;
     out254            :out std_logic;
     out255            :out std_logic;
     out256            :out std_logic;
     out257            :out std_logic;
     out258            :out std_logic;
     out259            :out std_logic;
     out260            :out std_logic;
     out261            :out std_logic;
     out262            :out std_logic;
     out263            :out std_logic;
     out264            :out std_logic;
     out265            :out std_logic;
     out266            :out std_logic;
     out267            :out std_logic;
     out268            :out std_logic;
     out269            :out std_logic;
     out270            :out std_logic;
     out271            :out std_logic;
     out272            :out std_logic;
     out273            :out std_logic;
     out274            :out std_logic;
     out275            :out std_logic;
     out276            :out std_logic;
     out277            :out std_logic;
     out278            :out std_logic;
     out279            :out std_logic;
     out280            :out std_logic;
     out281            :out std_logic;
     out282            :out std_logic;
     out283            :out std_logic;
     out284            :out std_logic;
     out285            :out std_logic;
     out286            :out std_logic;
     out287            :out std_logic;
     out288            :out std_logic;
     out289            :out std_logic;
     out290            :out std_logic;
     out291            :out std_logic;
     out292            :out std_logic;
     out293            :out std_logic;
     out294            :out std_logic;
     out295            :out std_logic;
     out296            :out std_logic;
     out297            :out std_logic;
     out298            :out std_logic;
     out299            :out std_logic;
     out300            :out std_logic;
     out301            :out std_logic;
     out302            :out std_logic;
     out303            :out std_logic;
     out304            :out std_logic;
     out305            :out std_logic;
     out306            :out std_logic;
     out307            :out std_logic;
     out308            :out std_logic;
     out309            :out std_logic;
     out310            :out std_logic;
     out311            :out std_logic;
     out312            :out std_logic;
     out313            :out std_logic;
     out314            :out std_logic;
     out315            :out std_logic;
     out316            :out std_logic;
     out317            :out std_logic;
     out318            :out std_logic;
     out319            :out std_logic;
     out320            :out std_logic;
     out321            :out std_logic;
     out322            :out std_logic;
     out323            :out std_logic;
     out324            :out std_logic;
     out325            :out std_logic;
     out326            :out std_logic;
     out327            :out std_logic;
     out328            :out std_logic;
     out329            :out std_logic;
     out330            :out std_logic;
     out331            :out std_logic;
     out332            :out std_logic;
     out333            :out std_logic;
     out334            :out std_logic;
     out335            :out std_logic;
     out336            :out std_logic;
     out337            :out std_logic;
     out338            :out std_logic;
     out339            :out std_logic;
     out340            :out std_logic;
     out341            :out std_logic;
     out342            :out std_logic;
     out343            :out std_logic;
     out344            :out std_logic;
     out345            :out std_logic;
     out346            :out std_logic;
     out347            :out std_logic;
     out348            :out std_logic;
     out349            :out std_logic;
     out350            :out std_logic;
     out351            :out std_logic;
     out352            :out std_logic;
     out353            :out std_logic;
     out354            :out std_logic;
     out355            :out std_logic;
     out356            :out std_logic;
     out357            :out std_logic;
     out358            :out std_logic;
     out359            :out std_logic;
     out360            :out std_logic;
     out361            :out std_logic;
     out362            :out std_logic;
     out363            :out std_logic;
     out364            :out std_logic;
     out365            :out std_logic;
     out366            :out std_logic;
     out367            :out std_logic;
     out368            :out std_logic;
     out369            :out std_logic;
     out370            :out std_logic;
     out371            :out std_logic;
     out372            :out std_logic;
     out373            :out std_logic;
     out374            :out std_logic;
     out375            :out std_logic;
     out376            :out std_logic;
     out377            :out std_logic;
     out378            :out std_logic;
     out379            :out std_logic;
     out380            :out std_logic;
     out381            :out std_logic;
     out382            :out std_logic;
     out383            :out std_logic;
     out384            :out std_logic;
     out385            :out std_logic;
     out386            :out std_logic;
     out387            :out std_logic;
     out388            :out std_logic;
     out389            :out std_logic;
     out390            :out std_logic;
     out391            :out std_logic;
     out392            :out std_logic;
     out393            :out std_logic;
     out394            :out std_logic;
     out395            :out std_logic;
     out396            :out std_logic;
     out397            :out std_logic;
     out398            :out std_logic;
     out399            :out std_logic;
     out400            :out std_logic;
     out401            :out std_logic;
     out402            :out std_logic;
     out403            :out std_logic;
     out404            :out std_logic;
     out405            :out std_logic;
     out406            :out std_logic;
     out407            :out std_logic;
     out408            :out std_logic;
     out409            :out std_logic;
     out410            :out std_logic;
     out411            :out std_logic;
     out412            :out std_logic;
     out413            :out std_logic;
     out414            :out std_logic;
     out415            :out std_logic;
     out416            :out std_logic;
     out417            :out std_logic;
     out418            :out std_logic;
     out419            :out std_logic;
     out420            :out std_logic;
     out421            :out std_logic;
     out422            :out std_logic;
     out423            :out std_logic;
     out424            :out std_logic;
     out425            :out std_logic;
     out426            :out std_logic;
     out427            :out std_logic;
     out428            :out std_logic;
     out429            :out std_logic;
     out430            :out std_logic;
     out431            :out std_logic;
     out432            :out std_logic;
     out433            :out std_logic;
     out434            :out std_logic;
     out435            :out std_logic;
     out436            :out std_logic;
     out437            :out std_logic;
     out438            :out std_logic;
     out439            :out std_logic;
     out440            :out std_logic;
     out441            :out std_logic;
     out442            :out std_logic;
     out443            :out std_logic;
     out444            :out std_logic;
     out445            :out std_logic;
     out446            :out std_logic;
     out447            :out std_logic;
     out448            :out std_logic;
     out449            :out std_logic;
     out450            :out std_logic;
     out451            :out std_logic;
     out452            :out std_logic;
     out453            :out std_logic;
     out454            :out std_logic;
     out455            :out std_logic;
     out456            :out std_logic;
     out457            :out std_logic;
     out458            :out std_logic;
     out459            :out std_logic;
     out460            :out std_logic;
     out461            :out std_logic;
     out462            :out std_logic;
     out463            :out std_logic;
     out464            :out std_logic;
     out465            :out std_logic;
     out466            :out std_logic;
     out467            :out std_logic;
     out468            :out std_logic;
     out469            :out std_logic;
     out470            :out std_logic;
     out471            :out std_logic;
     out472            :out std_logic;
     out473            :out std_logic;
     out474            :out std_logic;
     out475            :out std_logic;
     out476            :out std_logic;
     out477            :out std_logic;
     out478            :out std_logic;
     out479            :out std_logic;
     out480            :out std_logic;
     out481            :out std_logic;
     out482            :out std_logic;
     out483            :out std_logic;
     out484            :out std_logic;
     out485            :out std_logic;
     out486            :out std_logic;
     out487            :out std_logic;
     out488            :out std_logic;
     out489            :out std_logic;
     out490            :out std_logic;
     out491            :out std_logic;
     out492            :out std_logic;
     out493            :out std_logic;
     out494            :out std_logic;
     out495            :out std_logic;
     out496            :out std_logic;
     out497            :out std_logic;
     out498            :out std_logic;
     out499            :out std_logic;
     out500            :out std_logic;
     out501            :out std_logic;
     out502            :out std_logic;
     out503            :out std_logic;
     out504            :out std_logic;
     out505            :out std_logic;
     out506            :out std_logic;
     out507            :out std_logic;
     out508            :out std_logic;
     out509            :out std_logic;
     out510            :out std_logic;
     out511            :out std_logic;
     out512            :out std_logic;
     out513            :out std_logic;
     out514            :out std_logic;
     out515            :out std_logic;
     out516            :out std_logic;
     out517            :out std_logic;
     out518            :out std_logic;
     out519            :out std_logic;
     out520            :out std_logic;
     out521            :out std_logic;
     out522            :out std_logic;
     out523            :out std_logic;
     out524            :out std_logic;
     out525            :out std_logic;
     out526            :out std_logic;
     out527            :out std_logic;
     out528            :out std_logic;
     out529            :out std_logic;
     out530            :out std_logic;
     out531            :out std_logic;
     out532            :out std_logic;
     out533            :out std_logic;
     out534            :out std_logic;
     out535            :out std_logic;
     out536            :out std_logic;
     out537            :out std_logic;
     out538            :out std_logic;
     out539            :out std_logic;
     out540            :out std_logic;
     out541            :out std_logic;
     out542            :out std_logic;
     out543            :out std_logic;
     out544            :out std_logic;
     out545            :out std_logic;
     out546            :out std_logic;
     out547            :out std_logic;
     out548            :out std_logic;
     out549            :out std_logic;
     out550            :out std_logic;
     out551            :out std_logic;
     out552            :out std_logic;
     out553            :out std_logic;
     out554            :out std_logic;
     out555            :out std_logic;
     out556            :out std_logic;
     out557            :out std_logic;
     out558            :out std_logic;
     out559            :out std_logic;
     out560            :out std_logic;
     out561            :out std_logic;
     out562            :out std_logic;
     out563            :out std_logic;
     out564            :out std_logic;
     out565            :out std_logic;
     out566            :out std_logic;
     out567            :out std_logic;
     out568            :out std_logic;
     out569            :out std_logic;
     out570            :out std_logic;
     out571            :out std_logic;
     out572            :out std_logic;
     out573            :out std_logic;
     out574            :out std_logic;
     out575            :out std_logic;
     out576            :out std_logic;
     out577            :out std_logic;
     out578            :out std_logic;
     out579            :out std_logic;
     out580            :out std_logic;
     out581            :out std_logic;
     out582            :out std_logic;
     out583            :out std_logic;
     out584            :out std_logic;
     out585            :out std_logic;
     out586            :out std_logic;
     out587            :out std_logic;
     out588            :out std_logic;
     out589            :out std_logic;
     out590            :out std_logic;
     out591            :out std_logic;
     out592            :out std_logic;
     out593            :out std_logic;
     out594            :out std_logic;
     out595            :out std_logic;
     out596            :out std_logic;
     out597            :out std_logic;
     out598            :out std_logic;
     out599            :out std_logic;
     out600            :out std_logic;
     out601            :out std_logic;
     out602            :out std_logic;
     out603            :out std_logic;
     out604            :out std_logic;
     out605            :out std_logic;
     out606            :out std_logic;
     out607            :out std_logic;
     out608            :out std_logic;
     out609            :out std_logic;
     out610            :out std_logic;
     out611            :out std_logic;
     out612            :out std_logic;
     out613            :out std_logic;
     out614            :out std_logic;
     out615            :out std_logic;
     out616            :out std_logic;
     out617            :out std_logic;
     out618            :out std_logic;
     out619            :out std_logic;
     out620            :out std_logic;
     out621            :out std_logic;
     out622            :out std_logic;
     out623            :out std_logic;
     out624            :out std_logic;
     out625            :out std_logic;
     out626            :out std_logic;
     out627            :out std_logic;
     out628            :out std_logic;
     out629            :out std_logic;
     out630            :out std_logic;
     out631            :out std_logic;
     out632            :out std_logic;
     out633            :out std_logic;
     out634            :out std_logic;
     out635            :out std_logic;
     out636            :out std_logic;
     out637            :out std_logic;
     out638            :out std_logic;
     out639            :out std_logic;
     out640            :out std_logic;
     out641            :out std_logic;
     out642            :out std_logic;
     out643            :out std_logic;
     out644            :out std_logic;
     out645            :out std_logic;
     out646            :out std_logic;
     out647            :out std_logic;
     out648            :out std_logic;
     out649            :out std_logic;
     out650            :out std_logic;
     out651            :out std_logic;
     out652            :out std_logic;
     out653            :out std_logic;
     out654            :out std_logic;
     out655            :out std_logic;
     out656            :out std_logic;
     out657            :out std_logic;
     out658            :out std_logic;
     out659            :out std_logic;
     out660            :out std_logic;
     out661            :out std_logic;
     out662            :out std_logic;
     out663            :out std_logic;
     out664            :out std_logic;
     out665            :out std_logic;
     out666            :out std_logic;
     out667            :out std_logic;
     out668            :out std_logic;
     out669            :out std_logic;
     out670            :out std_logic;
     out671            :out std_logic;
     out672            :out std_logic;
     out673            :out std_logic;
     out674            :out std_logic;
     out675            :out std_logic;
     out676            :out std_logic;
     out677            :out std_logic;
     out678            :out std_logic;
     out679            :out std_logic;
     out680            :out std_logic;
     out681            :out std_logic;
     out682            :out std_logic;
     out683            :out std_logic;
     out684            :out std_logic;
     out685            :out std_logic;
     out686            :out std_logic;
     out687            :out std_logic;
     out688            :out std_logic;
     out689            :out std_logic;
     out690            :out std_logic;
     out691            :out std_logic;
     out692            :out std_logic;
     out693            :out std_logic;
     out694            :out std_logic;
     out695            :out std_logic;
     out696            :out std_logic;
     out697            :out std_logic;
     out698            :out std_logic;
     out699            :out std_logic;
     out700            :out std_logic;
     out701            :out std_logic;
     out702            :out std_logic;
     out703            :out std_logic;
     out704            :out std_logic;
     out705            :out std_logic;
     out706            :out std_logic;
     out707            :out std_logic;
     out708            :out std_logic;
     out709            :out std_logic;
     out710            :out std_logic;
     out711            :out std_logic;
     out712            :out std_logic;
     out713            :out std_logic;
     out714            :out std_logic;
     out715            :out std_logic;
     out716            :out std_logic;
     out717            :out std_logic;
     out718            :out std_logic;
     out719            :out std_logic;
     out720            :out std_logic;
     out721            :out std_logic;
     out722            :out std_logic;
     out723            :out std_logic;
     out724            :out std_logic;
     out725            :out std_logic;
     out726            :out std_logic;
     out727            :out std_logic;
     out728            :out std_logic;
     out729            :out std_logic;
     out730            :out std_logic;
     out731            :out std_logic;
     out732            :out std_logic;
     out733            :out std_logic;
     out734            :out std_logic;
     out735            :out std_logic;
     out736            :out std_logic;
     out737            :out std_logic;
     out738            :out std_logic;
     out739            :out std_logic;
     out740            :out std_logic;
     out741            :out std_logic;
     out742            :out std_logic;
     out743            :out std_logic;
     out744            :out std_logic;
     out745            :out std_logic;
     out746            :out std_logic;
     out747            :out std_logic;
     out748            :out std_logic;
     out749            :out std_logic;
     out750            :out std_logic;
     out751            :out std_logic;
     out752            :out std_logic;
     out753            :out std_logic;
     out754            :out std_logic;
     out755            :out std_logic;
     out756            :out std_logic;
     out757            :out std_logic;
     out758            :out std_logic;
     out759            :out std_logic;
     out760            :out std_logic;
     out761            :out std_logic;
     out762            :out std_logic;
     out763            :out std_logic;
     out764            :out std_logic;
     out765            :out std_logic;
     out766            :out std_logic;
     out767            :out std_logic;
     out768            :out std_logic;
     out769            :out std_logic;
     out770            :out std_logic;
     out771            :out std_logic;
     out772            :out std_logic;
     out773            :out std_logic;
     out774            :out std_logic;
     out775            :out std_logic;
     out776            :out std_logic;
     out777            :out std_logic;
     out778            :out std_logic;
     out779            :out std_logic;
     out780            :out std_logic;
     out781            :out std_logic;
     out782            :out std_logic;
     out783            :out std_logic;
     out784            :out std_logic;
     out785            :out std_logic;
     out786            :out std_logic;
     out787            :out std_logic;
     out788            :out std_logic;
     out789            :out std_logic;
     out790            :out std_logic;
     out791            :out std_logic;
     out792            :out std_logic;
     out793            :out std_logic;
     out794            :out std_logic;
     out795            :out std_logic;
     out796            :out std_logic;
     out797            :out std_logic;
     out798            :out std_logic;
     out799            :out std_logic;
     out800            :out std_logic;
     out801            :out std_logic;
     out802            :out std_logic;
     out803            :out std_logic;
     out804            :out std_logic;
     out805            :out std_logic;
     out806            :out std_logic;
     out807            :out std_logic;
     out808            :out std_logic;
     out809            :out std_logic;
     out810            :out std_logic;
     out811            :out std_logic;
     out812            :out std_logic;
     out813            :out std_logic;
     out814            :out std_logic;
     out815            :out std_logic;
     out816            :out std_logic;
     out817            :out std_logic;
     out818            :out std_logic;
     out819            :out std_logic;
     out820            :out std_logic;
     out821            :out std_logic;
     out822            :out std_logic;
     out823            :out std_logic;
     out824            :out std_logic;
     out825            :out std_logic;
     out826            :out std_logic;
     out827            :out std_logic;
     out828            :out std_logic;
     out829            :out std_logic;
     out830            :out std_logic;
     out831            :out std_logic;
     out832            :out std_logic;
     out833            :out std_logic;
     out834            :out std_logic;
     out835            :out std_logic;
     out836            :out std_logic;
     out837            :out std_logic;
     out838            :out std_logic;
     out839            :out std_logic;
     out840            :out std_logic;
     out841            :out std_logic;
     out842            :out std_logic;
     out843            :out std_logic;
     out844            :out std_logic;
     out845            :out std_logic;
     out846            :out std_logic;
     out847            :out std_logic;
     out848            :out std_logic;
     out849            :out std_logic;
     out850            :out std_logic;
     out851            :out std_logic;
     out852            :out std_logic;
     out853            :out std_logic;
     out854            :out std_logic;
     out855            :out std_logic;
     out856            :out std_logic;
     out857            :out std_logic;
     out858            :out std_logic;
     out859            :out std_logic;
     out860            :out std_logic;
     out861            :out std_logic;
     out862            :out std_logic;
     out863            :out std_logic;
     out864            :out std_logic;
     out865            :out std_logic;
     out866            :out std_logic;
     out867            :out std_logic;
     out868            :out std_logic;
     out869            :out std_logic;
     out870            :out std_logic;
     out871            :out std_logic;
     out872            :out std_logic;
     out873            :out std_logic;
     out874            :out std_logic;
     out875            :out std_logic;
     out876            :out std_logic;
     out877            :out std_logic;
     out878            :out std_logic;
     out879            :out std_logic;
     out880            :out std_logic;
     out881            :out std_logic;
     out882            :out std_logic;
     out883            :out std_logic;
     out884            :out std_logic;
     out885            :out std_logic;
     out886            :out std_logic;
     out887            :out std_logic;
     out888            :out std_logic;
     out889            :out std_logic;
     out890            :out std_logic;
     out891            :out std_logic;
     out892            :out std_logic;
     out893            :out std_logic;
     out894            :out std_logic;
     out895            :out std_logic;
     out896            :out std_logic;
     out897            :out std_logic;
     out898            :out std_logic;
     out899            :out std_logic;
     out900            :out std_logic;
     out901            :out std_logic;
     out902            :out std_logic;
     out903            :out std_logic;
     out904            :out std_logic;
     out905            :out std_logic;
     out906            :out std_logic;
     out907            :out std_logic;
     out908            :out std_logic;
     out909            :out std_logic;
     out910            :out std_logic;
     out911            :out std_logic;
     out912            :out std_logic;
     out913            :out std_logic;
     out914            :out std_logic;
     out915            :out std_logic;
     out916            :out std_logic;
     out917            :out std_logic;
     out918            :out std_logic;
     out919            :out std_logic;
     out920            :out std_logic;
     out921            :out std_logic;
     out922            :out std_logic;
     out923            :out std_logic;
     out924            :out std_logic;
     out925            :out std_logic;
     out926            :out std_logic;
     out927            :out std_logic;
     out928            :out std_logic;
     out929            :out std_logic;
     out930            :out std_logic;
     out931            :out std_logic;
     out932            :out std_logic;
     out933            :out std_logic;
     out934            :out std_logic;
     out935            :out std_logic;
     out936            :out std_logic;
     out937            :out std_logic;
     out938            :out std_logic;
     out939            :out std_logic;
     out940            :out std_logic;
     out941            :out std_logic;
     out942            :out std_logic;
     out943            :out std_logic;
     out944            :out std_logic;
     out945            :out std_logic;
     out946            :out std_logic;
     out947            :out std_logic;
     out948            :out std_logic;
     out949            :out std_logic;
     out950            :out std_logic;
     out951            :out std_logic;
     out952            :out std_logic;
     out953            :out std_logic;
     out954            :out std_logic;
     out955            :out std_logic;
     out956            :out std_logic;
     out957            :out std_logic;
     out958            :out std_logic;
     out959            :out std_logic;
     out960            :out std_logic;
     out961            :out std_logic;
     out962            :out std_logic;
     out963            :out std_logic;
     out964            :out std_logic;
     out965            :out std_logic;
     out966            :out std_logic;
     out967            :out std_logic;
     out968            :out std_logic;
     out969            :out std_logic;
     out970            :out std_logic;
     out971            :out std_logic;
     out972            :out std_logic;
     out973            :out std_logic;
     out974            :out std_logic;
     out975            :out std_logic;
     out976            :out std_logic;
     out977            :out std_logic;
     out978            :out std_logic;
     out979            :out std_logic;
     out980            :out std_logic;
     out981            :out std_logic;
     out982            :out std_logic;
     out983            :out std_logic;
     out984            :out std_logic;
     out985            :out std_logic;
     out986            :out std_logic;
     out987            :out std_logic;
     out988            :out std_logic;
     out989            :out std_logic;
     out990            :out std_logic;
     out991            :out std_logic;
     out992            :out std_logic;
     out993            :out std_logic;
     out994            :out std_logic;
     out995            :out std_logic;
     out996            :out std_logic;
     out997            :out std_logic;
     out998            :out std_logic;
     out999            :out std_logic;
     out1000            :out std_logic;
     out1001            :out std_logic;
     out1002            :out std_logic;
     out1003            :out std_logic;
     out1004            :out std_logic;
     out1005            :out std_logic;
     out1006            :out std_logic;
     out1007            :out std_logic;
     out1008            :out std_logic;
     out1009            :out std_logic;
     out1010            :out std_logic;
     out1011            :out std_logic;
     out1012            :out std_logic;
     out1013            :out std_logic;
     out1014            :out std_logic;
     out1015            :out std_logic;
     out1016            :out std_logic;
     out1017            :out std_logic;
     out1018            :out std_logic;
     out1019            :out std_logic;
     out1020            :out std_logic;
     out1021            :out std_logic;
     out1022            :out std_logic;
     out1023            :out std_logic;
     out1024            :out std_logic;
     out1025            :out std_logic;
     out1026            :out std_logic;
     out1027            :out std_logic;
     out1028            :out std_logic;
     out1029            :out std_logic;
     out1030            :out std_logic;
     out1031            :out std_logic;
     out1032            :out std_logic;
     out1033            :out std_logic;
     out1034            :out std_logic;
     out1035            :out std_logic;
     out1036            :out std_logic;
     out1037            :out std_logic;
     out1038            :out std_logic;
     out1039            :out std_logic;
     out1040            :out std_logic;
     out1041            :out std_logic;
     out1042            :out std_logic;
     out1043            :out std_logic;
     out1044            :out std_logic;
     out1045            :out std_logic;
     out1046            :out std_logic;
     out1047            :out std_logic;
     out1048            :out std_logic;
     out1049            :out std_logic;
     out1050            :out std_logic;
     out1051            :out std_logic;
     out1052            :out std_logic;
     out1053            :out std_logic;
     out1054            :out std_logic;
     out1055            :out std_logic;
     out1056            :out std_logic;
     out1057            :out std_logic;
     out1058            :out std_logic;
     out1059            :out std_logic;
     out1060            :out std_logic;
     out1061            :out std_logic;
     out1062            :out std_logic;
     out1063            :out std_logic;
     out1064            :out std_logic;
     out1065            :out std_logic;
     out1066            :out std_logic;
     out1067            :out std_logic;
     out1068            :out std_logic;
     out1069            :out std_logic;
     out1070            :out std_logic;
     out1071            :out std_logic;
     out1072            :out std_logic;
     out1073            :out std_logic;
     out1074            :out std_logic;
     out1075            :out std_logic;
     out1076            :out std_logic;
     out1077            :out std_logic;
     out1078            :out std_logic;
     out1079            :out std_logic;
     out1080            :out std_logic;
     out1081            :out std_logic;
     out1082            :out std_logic;
     out1083            :out std_logic;
     out1084            :out std_logic;
     out1085            :out std_logic;
     out1086            :out std_logic;
     out1087            :out std_logic;
     out1088            :out std_logic;
     out1089            :out std_logic;
     out1090            :out std_logic;
     out1091            :out std_logic;
     out1092            :out std_logic;
     out1093            :out std_logic;
     out1094            :out std_logic;
     out1095            :out std_logic;
     out1096            :out std_logic;
     out1097            :out std_logic;
     out1098            :out std_logic;
     out1099            :out std_logic;
     out1100            :out std_logic;
     out1101            :out std_logic;
     out1102            :out std_logic;
     out1103            :out std_logic;
     out1104            :out std_logic;
     out1105            :out std_logic;
     out1106            :out std_logic;
     out1107            :out std_logic;
     out1108            :out std_logic;
     out1109            :out std_logic;
     out1110            :out std_logic;
     out1111            :out std_logic;
     out1112            :out std_logic;
     out1113            :out std_logic;
     out1114            :out std_logic;
     out1115            :out std_logic;
     out1116            :out std_logic;
     out1117            :out std_logic;
     out1118            :out std_logic;
     out1119            :out std_logic;
     out1120            :out std_logic;
     out1121            :out std_logic;
     out1122            :out std_logic;
     out1123            :out std_logic;
     out1124            :out std_logic;
     out1125            :out std_logic;
     out1126            :out std_logic;
     out1127            :out std_logic;
     out1128            :out std_logic;
     out1129            :out std_logic;
     out1130            :out std_logic;
     out1131            :out std_logic;
     out1132            :out std_logic;
     out1133            :out std_logic;
     out1134            :out std_logic;
     out1135            :out std_logic;
     out1136            :out std_logic;
     out1137            :out std_logic;
     out1138            :out std_logic;
     out1139            :out std_logic;
     out1140            :out std_logic;
     out1141            :out std_logic;
     out1142            :out std_logic;
     out1143            :out std_logic;
     out1144            :out std_logic;
     out1145            :out std_logic;
     out1146            :out std_logic;
     out1147            :out std_logic;
     out1148            :out std_logic;
     out1149            :out std_logic;
     out1150            :out std_logic;
     out1151            :out std_logic;
     out1152            :out std_logic;
     out1153            :out std_logic;
     out1154            :out std_logic;
     out1155            :out std_logic;
     out1156            :out std_logic;
     out1157            :out std_logic;
     out1158            :out std_logic;
     out1159            :out std_logic;
     out1160            :out std_logic;
     out1161            :out std_logic;
     out1162            :out std_logic;
     out1163            :out std_logic;
     out1164            :out std_logic;
     out1165            :out std_logic;
     out1166            :out std_logic;
     out1167            :out std_logic;
     out1168            :out std_logic;
     out1169            :out std_logic;
     out1170            :out std_logic;
     out1171            :out std_logic;
     out1172            :out std_logic;
     out1173            :out std_logic;
     out1174            :out std_logic;
     out1175            :out std_logic;
     out1176            :out std_logic;
     out1177            :out std_logic;
     out1178            :out std_logic;
     out1179            :out std_logic;
     out1180            :out std_logic;
     out1181            :out std_logic;
     out1182            :out std_logic;
     out1183            :out std_logic;
     out1184            :out std_logic;
     out1185            :out std_logic;
     out1186            :out std_logic;
     out1187            :out std_logic;
     out1188            :out std_logic;
     out1189            :out std_logic;
     out1190            :out std_logic;
     out1191            :out std_logic;
     out1192            :out std_logic;
     out1193            :out std_logic;
     out1194            :out std_logic;
     out1195            :out std_logic;
     out1196            :out std_logic;
     out1197            :out std_logic;
     out1198            :out std_logic;
     out1199            :out std_logic;
     out1200            :out std_logic;
     out1201            :out std_logic;
     out1202            :out std_logic;
     out1203            :out std_logic;
     out1204            :out std_logic;
     out1205            :out std_logic;
     out1206            :out std_logic;
     out1207            :out std_logic;
     out1208            :out std_logic;
     out1209            :out std_logic;
     out1210            :out std_logic;
     out1211            :out std_logic;
     out1212            :out std_logic;
     out1213            :out std_logic;
     out1214            :out std_logic;
     out1215            :out std_logic;
     out1216            :out std_logic;
     out1217            :out std_logic;
     out1218            :out std_logic;
     out1219            :out std_logic;
     out1220            :out std_logic;
     out1221            :out std_logic;
     out1222            :out std_logic;
     out1223            :out std_logic;
     out1224            :out std_logic;
     out1225            :out std_logic;
     out1226            :out std_logic;
     out1227            :out std_logic;
     out1228            :out std_logic;
     out1229            :out std_logic;
     out1230            :out std_logic;
     out1231            :out std_logic;
     out1232            :out std_logic;
     out1233            :out std_logic;
     out1234            :out std_logic;
     out1235            :out std_logic;
     out1236            :out std_logic;
     out1237            :out std_logic;
     out1238            :out std_logic;
     out1239            :out std_logic;
     out1240            :out std_logic;
     out1241            :out std_logic;
     out1242            :out std_logic;
     out1243            :out std_logic;
     out1244            :out std_logic;
     out1245            :out std_logic;
     out1246            :out std_logic;
     out1247            :out std_logic;
     out1248            :out std_logic;
     out1249            :out std_logic;
     out1250            :out std_logic;
     out1251            :out std_logic;
     out1252            :out std_logic;
     out1253            :out std_logic;
     out1254            :out std_logic;
     out1255            :out std_logic;
     out1256            :out std_logic;
     out1257            :out std_logic;
     out1258            :out std_logic;
     out1259            :out std_logic;
     out1260            :out std_logic;
     out1261            :out std_logic;
     out1262            :out std_logic;
     out1263            :out std_logic;
     out1264            :out std_logic;
     out1265            :out std_logic;
     out1266            :out std_logic;
     out1267            :out std_logic;
     out1268            :out std_logic;
     out1269            :out std_logic;
     out1270            :out std_logic;
     out1271            :out std_logic;
     out1272            :out std_logic;
     out1273            :out std_logic;
     out1274            :out std_logic;
     out1275            :out std_logic;
     out1276            :out std_logic;
     out1277            :out std_logic;
     out1278            :out std_logic;
     out1279            :out std_logic;
     out1280            :out std_logic;
     out1281            :out std_logic;
     out1282            :out std_logic;
     out1283            :out std_logic;
     out1284            :out std_logic;
     out1285            :out std_logic;
     out1286            :out std_logic;
     out1287            :out std_logic;
     out1288            :out std_logic;
     out1289            :out std_logic;
     out1290            :out std_logic;
     out1291            :out std_logic;
     out1292            :out std_logic;
     out1293            :out std_logic;
     out1294            :out std_logic;
     out1295            :out std_logic;
     out1296            :out std_logic;
     out1297            :out std_logic;
     out1298            :out std_logic;
     out1299            :out std_logic;
     out1300            :out std_logic;
     out1301            :out std_logic;
     out1302            :out std_logic;
     out1303            :out std_logic;
     out1304            :out std_logic;
     out1305            :out std_logic;
     out1306            :out std_logic;
     out1307            :out std_logic;
     out1308            :out std_logic;
     out1309            :out std_logic;
     out1310            :out std_logic;
     out1311            :out std_logic;
     out1312            :out std_logic;
     out1313            :out std_logic;
     out1314            :out std_logic;
     out1315            :out std_logic;
     out1316            :out std_logic;
     out1317            :out std_logic;
     out1318            :out std_logic;
     out1319            :out std_logic;
     out1320            :out std_logic;
     out1321            :out std_logic;
     out1322            :out std_logic;
     out1323            :out std_logic;
     out1324            :out std_logic;
     out1325            :out std_logic;
     out1326            :out std_logic;
     out1327            :out std_logic;
     out1328            :out std_logic;
     out1329            :out std_logic;
     out1330            :out std_logic;
     out1331            :out std_logic;
     out1332            :out std_logic;
     out1333            :out std_logic;
     out1334            :out std_logic;
     out1335            :out std_logic;
     out1336            :out std_logic;
     out1337            :out std_logic;
     out1338            :out std_logic;
     out1339            :out std_logic;
     out1340            :out std_logic;
     out1341            :out std_logic;
     out1342            :out std_logic;
     out1343            :out std_logic;
     out1344            :out std_logic;
     out1345            :out std_logic;
     out1346            :out std_logic;
     out1347            :out std_logic;
     out1348            :out std_logic;
     out1349            :out std_logic;
     out1350            :out std_logic;
     out1351            :out std_logic;
     out1352            :out std_logic;
     out1353            :out std_logic;
     out1354            :out std_logic;
     out1355            :out std_logic;
     out1356            :out std_logic;
     out1357            :out std_logic;
     out1358            :out std_logic;
     out1359            :out std_logic;
     out1360            :out std_logic;
     out1361            :out std_logic;
     out1362            :out std_logic;
     out1363            :out std_logic;
     out1364            :out std_logic;
     out1365            :out std_logic;
     out1366            :out std_logic;
     out1367            :out std_logic;
     out1368            :out std_logic;
     out1369            :out std_logic;
     out1370            :out std_logic;
     out1371            :out std_logic;
     out1372            :out std_logic;
     out1373            :out std_logic;
     out1374            :out std_logic;
     out1375            :out std_logic;
     out1376            :out std_logic;
     out1377            :out std_logic;
     out1378            :out std_logic;
     out1379            :out std_logic;
     out1380            :out std_logic;
     out1381            :out std_logic;
     out1382            :out std_logic;
     out1383            :out std_logic;
     out1384            :out std_logic;
     out1385            :out std_logic;
     out1386            :out std_logic;
     out1387            :out std_logic;
     out1388            :out std_logic;
     out1389            :out std_logic;
     out1390            :out std_logic;
     out1391            :out std_logic;
     out1392            :out std_logic;
     out1393            :out std_logic;
     out1394            :out std_logic;
     out1395            :out std_logic;
     out1396            :out std_logic;
     out1397            :out std_logic;
     out1398            :out std_logic;
     out1399            :out std_logic;
     out1400            :out std_logic;
     out1401            :out std_logic;
     out1402            :out std_logic;
     out1403            :out std_logic;
     out1404            :out std_logic;
     out1405            :out std_logic;
     out1406            :out std_logic;
     out1407            :out std_logic;
     out1408            :out std_logic;
     out1409            :out std_logic;
     out1410            :out std_logic;
     out1411            :out std_logic;
     out1412            :out std_logic;
     out1413            :out std_logic;
     out1414            :out std_logic;
     out1415            :out std_logic;
     out1416            :out std_logic;
     out1417            :out std_logic;
     out1418            :out std_logic;
     out1419            :out std_logic;
     out1420            :out std_logic;
     out1421            :out std_logic;
     out1422            :out std_logic;
     out1423            :out std_logic;
     out1424            :out std_logic;
     out1425            :out std_logic;
     out1426            :out std_logic;
     out1427            :out std_logic;
     out1428            :out std_logic;
     out1429            :out std_logic;
     out1430            :out std_logic;
     out1431            :out std_logic;
     out1432            :out std_logic;
     out1433            :out std_logic;
     out1434            :out std_logic;
     out1435            :out std_logic;
     out1436            :out std_logic;
     out1437            :out std_logic;
     out1438            :out std_logic;
     out1439            :out std_logic;
     out1440            :out std_logic;
     out1441            :out std_logic;
     out1442            :out std_logic;
     out1443            :out std_logic;
     out1444            :out std_logic;
     out1445            :out std_logic;
     out1446            :out std_logic;
     out1447            :out std_logic;
     out1448            :out std_logic;
     out1449            :out std_logic;
     out1450            :out std_logic;
     out1451            :out std_logic;
     out1452            :out std_logic;
     out1453            :out std_logic;
     out1454            :out std_logic;
     out1455            :out std_logic;
     out1456            :out std_logic;
     out1457            :out std_logic;
     out1458            :out std_logic;
     out1459            :out std_logic;
     out1460            :out std_logic;
     out1461            :out std_logic;
     out1462            :out std_logic;
     out1463            :out std_logic;
     out1464            :out std_logic;
     out1465            :out std_logic;
     out1466            :out std_logic;
     out1467            :out std_logic;
     out1468            :out std_logic;
     out1469            :out std_logic;
     out1470            :out std_logic;
     out1471            :out std_logic;
     out1472            :out std_logic;
     out1473            :out std_logic;
     out1474            :out std_logic;
     out1475            :out std_logic;
     out1476            :out std_logic;
     out1477            :out std_logic;
     out1478            :out std_logic;
     out1479            :out std_logic;
     out1480            :out std_logic;
     out1481            :out std_logic;
     out1482            :out std_logic;
     out1483            :out std_logic;
     out1484            :out std_logic;
     out1485            :out std_logic;
     out1486            :out std_logic;
     out1487            :out std_logic;
     out1488            :out std_logic;
     out1489            :out std_logic;
     out1490            :out std_logic;
     out1491            :out std_logic;
     out1492            :out std_logic;
     out1493            :out std_logic;
     out1494            :out std_logic;
     out1495            :out std_logic;
     out1496            :out std_logic;
     out1497            :out std_logic;
     out1498            :out std_logic;
     out1499            :out std_logic;
     out1500            :out std_logic;
     out1501            :out std_logic;
     out1502            :out std_logic;
     out1503            :out std_logic;
     out1504            :out std_logic;
     out1505            :out std_logic;
     out1506            :out std_logic;
     out1507            :out std_logic;
     out1508            :out std_logic;
     out1509            :out std_logic;
     out1510            :out std_logic;
     out1511            :out std_logic;
     out1512            :out std_logic;
     out1513            :out std_logic;
     out1514            :out std_logic;
     out1515            :out std_logic;
     out1516            :out std_logic;
     out1517            :out std_logic;
     out1518            :out std_logic;
     out1519            :out std_logic;
     out1520            :out std_logic;
     out1521            :out std_logic;
     out1522            :out std_logic;
     out1523            :out std_logic;
     out1524            :out std_logic;
     out1525            :out std_logic;
     out1526            :out std_logic;
     out1527            :out std_logic;
     out1528            :out std_logic;
     out1529            :out std_logic;
     out1530            :out std_logic;
     out1531            :out std_logic;
     out1532            :out std_logic;
     out1533            :out std_logic;
     out1534            :out std_logic;
     out1535            :out std_logic;
     out1536            :out std_logic;
     out1537            :out std_logic;
     out1538            :out std_logic;
     out1539            :out std_logic;
     out1540            :out std_logic;
     out1541            :out std_logic;
     out1542            :out std_logic;
     out1543            :out std_logic;
     out1544            :out std_logic;
     out1545            :out std_logic;
     out1546            :out std_logic;
     out1547            :out std_logic;
     out1548            :out std_logic;
     out1549            :out std_logic;
     out1550            :out std_logic;
     out1551            :out std_logic;
     out1552            :out std_logic;
     out1553            :out std_logic;
     out1554            :out std_logic;
     out1555            :out std_logic;
     out1556            :out std_logic;
     out1557            :out std_logic;
     out1558            :out std_logic;
     out1559            :out std_logic;
     out1560            :out std_logic;
     out1561            :out std_logic;
     out1562            :out std_logic;
     out1563            :out std_logic;
     out1564            :out std_logic;
     out1565            :out std_logic;
     out1566            :out std_logic;
     out1567            :out std_logic;
     out1568            :out std_logic;
     out1569            :out std_logic;
     out1570            :out std_logic;
     out1571            :out std_logic;
     out1572            :out std_logic;
     out1573            :out std_logic;
     out1574            :out std_logic;
     out1575            :out std_logic;
     out1576            :out std_logic;
     out1577            :out std_logic;
     out1578            :out std_logic;
     out1579            :out std_logic;
     out1580            :out std_logic;
     out1581            :out std_logic;
     out1582            :out std_logic;
     out1583            :out std_logic;
     out1584            :out std_logic;
     out1585            :out std_logic;
     out1586            :out std_logic;
     out1587            :out std_logic;
     out1588            :out std_logic;
     out1589            :out std_logic;
     out1590            :out std_logic;
     out1591            :out std_logic;
     out1592            :out std_logic;
     out1593            :out std_logic;
     out1594            :out std_logic;
     out1595            :out std_logic;
     out1596            :out std_logic;
     out1597            :out std_logic;
     out1598            :out std_logic;
     out1599            :out std_logic;
     out1600            :out std_logic;
     out1601            :out std_logic;
     out1602            :out std_logic;
     out1603            :out std_logic;
     out1604            :out std_logic;
     out1605            :out std_logic;
     out1606            :out std_logic;
     out1607            :out std_logic;
     out1608            :out std_logic;
     out1609            :out std_logic;
     out1610            :out std_logic;
     out1611            :out std_logic;
     out1612            :out std_logic;
     out1613            :out std_logic;
     out1614            :out std_logic;
     out1615            :out std_logic;
     out1616            :out std_logic;
     out1617            :out std_logic;
     out1618            :out std_logic;
     out1619            :out std_logic;
     out1620            :out std_logic;
     out1621            :out std_logic;
     out1622            :out std_logic;
     out1623            :out std_logic;
     out1624            :out std_logic;
     out1625            :out std_logic;
     out1626            :out std_logic;
     out1627            :out std_logic;
     out1628            :out std_logic;
     out1629            :out std_logic;
     out1630            :out std_logic;
     out1631            :out std_logic;
     out1632            :out std_logic;
     out1633            :out std_logic;
     out1634            :out std_logic;
     out1635            :out std_logic;
     out1636            :out std_logic;
     out1637            :out std_logic;
     out1638            :out std_logic;
     out1639            :out std_logic;
     out1640            :out std_logic;
     out1641            :out std_logic;
     out1642            :out std_logic;
     out1643            :out std_logic;
     out1644            :out std_logic;
     out1645            :out std_logic;
     out1646            :out std_logic;
     out1647            :out std_logic;
     out1648            :out std_logic;
     out1649            :out std_logic;
     out1650            :out std_logic;
     out1651            :out std_logic;
     out1652            :out std_logic;
     out1653            :out std_logic;
     out1654            :out std_logic;
     out1655            :out std_logic;
     out1656            :out std_logic;
     out1657            :out std_logic;
     out1658            :out std_logic;
     out1659            :out std_logic;
     out1660            :out std_logic;
     out1661            :out std_logic;
     out1662            :out std_logic;
     out1663            :out std_logic;
     out1664            :out std_logic;
     out1665            :out std_logic;
     out1666            :out std_logic;
     out1667            :out std_logic;
     out1668            :out std_logic;
     out1669            :out std_logic;
     out1670            :out std_logic;
     out1671            :out std_logic;
     out1672            :out std_logic;
     out1673            :out std_logic;
     out1674            :out std_logic;
     out1675            :out std_logic;
     out1676            :out std_logic;
     out1677            :out std_logic;
     out1678            :out std_logic;
     out1679            :out std_logic;
     out1680            :out std_logic;
     out1681            :out std_logic;
     out1682            :out std_logic;
     out1683            :out std_logic;
     out1684            :out std_logic;
     out1685            :out std_logic;
     out1686            :out std_logic;
     out1687            :out std_logic;
     out1688            :out std_logic;
     out1689            :out std_logic;
     out1690            :out std_logic;
     out1691            :out std_logic;
     out1692            :out std_logic;
     out1693            :out std_logic;
     out1694            :out std_logic;
     out1695            :out std_logic;
     out1696            :out std_logic;
     out1697            :out std_logic;
     out1698            :out std_logic;
     out1699            :out std_logic;
     out1700            :out std_logic;
     out1701            :out std_logic;
     out1702            :out std_logic;
     out1703            :out std_logic;
     out1704            :out std_logic;
     out1705            :out std_logic;
     out1706            :out std_logic;
     out1707            :out std_logic;
     out1708            :out std_logic;
     out1709            :out std_logic;
     out1710            :out std_logic;
     out1711            :out std_logic;
     out1712            :out std_logic;
     out1713            :out std_logic;
     out1714            :out std_logic;
     out1715            :out std_logic;
     out1716            :out std_logic;
     out1717            :out std_logic;
     out1718            :out std_logic;
     out1719            :out std_logic;
     out1720            :out std_logic;
     out1721            :out std_logic;
     out1722            :out std_logic;
     out1723            :out std_logic;
     out1724            :out std_logic;
     out1725            :out std_logic;
     out1726            :out std_logic;
     out1727            :out std_logic;
     out1728            :out std_logic;
     out1729            :out std_logic;
     out1730            :out std_logic;
     out1731            :out std_logic;
     out1732            :out std_logic;
     out1733            :out std_logic;
     out1734            :out std_logic;
     out1735            :out std_logic;
     out1736            :out std_logic;
     out1737            :out std_logic;
     out1738            :out std_logic;
     out1739            :out std_logic;
     out1740            :out std_logic;
     out1741            :out std_logic;
     out1742            :out std_logic;
     out1743            :out std_logic;
     out1744            :out std_logic;
     out1745            :out std_logic;
     out1746            :out std_logic;
     out1747            :out std_logic;
     out1748            :out std_logic;
     out1749            :out std_logic;
     out1750            :out std_logic;
     out1751            :out std_logic;
     out1752            :out std_logic;
     out1753            :out std_logic;
     out1754            :out std_logic;
     out1755            :out std_logic;
     out1756            :out std_logic;
     out1757            :out std_logic;
     out1758            :out std_logic;
     out1759            :out std_logic;
     out1760            :out std_logic;
     out1761            :out std_logic;
     out1762            :out std_logic;
     out1763            :out std_logic;
     out1764            :out std_logic;
     out1765            :out std_logic;
     out1766            :out std_logic;
     out1767            :out std_logic;
     out1768            :out std_logic;
     out1769            :out std_logic;
     out1770            :out std_logic;
     out1771            :out std_logic;
     out1772            :out std_logic;
     out1773            :out std_logic;
     out1774            :out std_logic;
     out1775            :out std_logic;
     out1776            :out std_logic;
     out1777            :out std_logic;
     out1778            :out std_logic;
     out1779            :out std_logic;
     out1780            :out std_logic;
     out1781            :out std_logic;
     out1782            :out std_logic;
     out1783            :out std_logic;
     out1784            :out std_logic;
     out1785            :out std_logic;
     out1786            :out std_logic;
     out1787            :out std_logic;
     out1788            :out std_logic;
     out1789            :out std_logic;
     out1790            :out std_logic;
     out1791            :out std_logic;
     out1792            :out std_logic;
     out1793            :out std_logic;
     out1794            :out std_logic;
     out1795            :out std_logic;
     out1796            :out std_logic;
     out1797            :out std_logic;
     out1798            :out std_logic;
     out1799            :out std_logic;
     out1800            :out std_logic;
     out1801            :out std_logic;
     out1802            :out std_logic;
     out1803            :out std_logic;
     out1804            :out std_logic;
     out1805            :out std_logic;
     out1806            :out std_logic;
     out1807            :out std_logic;
     out1808            :out std_logic;
     out1809            :out std_logic;
     out1810            :out std_logic;
     out1811            :out std_logic;
     out1812            :out std_logic;
     out1813            :out std_logic;
     out1814            :out std_logic;
     out1815            :out std_logic;
     out1816            :out std_logic;
     out1817            :out std_logic;
     out1818            :out std_logic;
     out1819            :out std_logic;
     out1820            :out std_logic;
     out1821            :out std_logic;
     out1822            :out std_logic;
     out1823            :out std_logic;
     out1824            :out std_logic;
     out1825            :out std_logic;
     out1826            :out std_logic;
     out1827            :out std_logic;
     out1828            :out std_logic;
     out1829            :out std_logic;
     out1830            :out std_logic;
     out1831            :out std_logic;
     out1832            :out std_logic;
     out1833            :out std_logic;
     out1834            :out std_logic;
     out1835            :out std_logic;
     out1836            :out std_logic;
     out1837            :out std_logic;
     out1838            :out std_logic;
     out1839            :out std_logic;
     out1840            :out std_logic;
     out1841            :out std_logic;
     out1842            :out std_logic;
     out1843            :out std_logic;
     out1844            :out std_logic;
     out1845            :out std_logic;
     out1846            :out std_logic;
     out1847            :out std_logic;
     out1848            :out std_logic;
     out1849            :out std_logic;
     out1850            :out std_logic;
     out1851            :out std_logic;
     out1852            :out std_logic;
     out1853            :out std_logic;
     out1854            :out std_logic;
     out1855            :out std_logic;
     out1856            :out std_logic;
     out1857            :out std_logic;
     out1858            :out std_logic;
     out1859            :out std_logic;
     out1860            :out std_logic;
     out1861            :out std_logic;
     out1862            :out std_logic;
     out1863            :out std_logic;
     out1864            :out std_logic;
     out1865            :out std_logic;
     out1866            :out std_logic;
     out1867            :out std_logic;
     out1868            :out std_logic;
     out1869            :out std_logic;
     out1870            :out std_logic;
     out1871            :out std_logic;
     out1872            :out std_logic;
     out1873            :out std_logic;
     out1874            :out std_logic;
     out1875            :out std_logic;
     out1876            :out std_logic;
     out1877            :out std_logic;
     out1878            :out std_logic;
     out1879            :out std_logic;
     out1880            :out std_logic;
     out1881            :out std_logic;
     out1882            :out std_logic;
     out1883            :out std_logic;
     out1884            :out std_logic;
     out1885            :out std_logic;
     out1886            :out std_logic;
     out1887            :out std_logic;
     out1888            :out std_logic;
     out1889            :out std_logic;
     out1890            :out std_logic;
     out1891            :out std_logic;
     out1892            :out std_logic;
     out1893            :out std_logic;
     out1894            :out std_logic;
     out1895            :out std_logic;
     out1896            :out std_logic;
     out1897            :out std_logic;
     out1898            :out std_logic;
     out1899            :out std_logic;
     out1900            :out std_logic;
     out1901            :out std_logic;
     out1902            :out std_logic;
     out1903            :out std_logic;
     out1904            :out std_logic;
     out1905            :out std_logic;
     out1906            :out std_logic;
     out1907            :out std_logic;
     out1908            :out std_logic;
     out1909            :out std_logic;
     out1910            :out std_logic;
     out1911            :out std_logic;
     out1912            :out std_logic;
     out1913            :out std_logic;
     out1914            :out std_logic;
     out1915            :out std_logic;
     out1916            :out std_logic;
     out1917            :out std_logic;
     out1918            :out std_logic;
     out1919            :out std_logic;
     out1920            :out std_logic;
     out1921            :out std_logic;
     out1922            :out std_logic;
     out1923            :out std_logic;
     out1924            :out std_logic;
     out1925            :out std_logic;
     out1926            :out std_logic;
     out1927            :out std_logic;
     out1928            :out std_logic;
     out1929            :out std_logic;
     out1930            :out std_logic;
     out1931            :out std_logic;
     out1932            :out std_logic;
     out1933            :out std_logic;
     out1934            :out std_logic;
     out1935            :out std_logic;
     out1936            :out std_logic;
     out1937            :out std_logic;
     out1938            :out std_logic;
     out1939            :out std_logic;
     out1940            :out std_logic;
     out1941            :out std_logic;
     out1942            :out std_logic;
     out1943            :out std_logic;
     out1944            :out std_logic;
     out1945            :out std_logic;
     out1946            :out std_logic;
     out1947            :out std_logic;
     out1948            :out std_logic;
     out1949            :out std_logic;
     out1950            :out std_logic;
     out1951            :out std_logic;
     out1952            :out std_logic;
     out1953            :out std_logic;
     out1954            :out std_logic;
     out1955            :out std_logic;
     out1956            :out std_logic;
     out1957            :out std_logic;
     out1958            :out std_logic;
     out1959            :out std_logic;
     out1960            :out std_logic;
     out1961            :out std_logic;
     out1962            :out std_logic;
     out1963            :out std_logic;
     out1964            :out std_logic;
     out1965            :out std_logic;
     out1966            :out std_logic;
     out1967            :out std_logic;
     out1968            :out std_logic;
     out1969            :out std_logic;
     out1970            :out std_logic;
     out1971            :out std_logic;
     out1972            :out std_logic;
     out1973            :out std_logic;
     out1974            :out std_logic;
     out1975            :out std_logic;
     out1976            :out std_logic;
     out1977            :out std_logic;
     out1978            :out std_logic;
     out1979            :out std_logic;
     out1980            :out std_logic;
     out1981            :out std_logic;
     out1982            :out std_logic;
     out1983            :out std_logic;
     out1984            :out std_logic;
     out1985            :out std_logic;
     out1986            :out std_logic;
     out1987            :out std_logic;
     out1988            :out std_logic;
     out1989            :out std_logic;
     out1990            :out std_logic;
     out1991            :out std_logic;
     out1992            :out std_logic;
     out1993            :out std_logic;
     out1994            :out std_logic;
     out1995            :out std_logic;
     out1996            :out std_logic;
     out1997            :out std_logic;
     out1998            :out std_logic;
     out1999            :out std_logic;
     out2000            :out std_logic;
     out2001            :out std_logic;
     out2002            :out std_logic;
     out2003            :out std_logic;
     out2004            :out std_logic;
     out2005            :out std_logic;
     out2006            :out std_logic;
     out2007            :out std_logic;
     out2008            :out std_logic;
     out2009            :out std_logic;
     out2010            :out std_logic;
     out2011            :out std_logic;
     out2012            :out std_logic;
     out2013            :out std_logic;
     out2014            :out std_logic;
     out2015            :out std_logic;
     out2016            :out std_logic;
     out2017            :out std_logic;
     out2018            :out std_logic;
     out2019            :out std_logic;
     out2020            :out std_logic;
     out2021            :out std_logic;
     out2022            :out std_logic;
     out2023            :out std_logic;
     out2024            :out std_logic;
     out2025            :out std_logic;
     out2026            :out std_logic;
     out2027            :out std_logic;
     out2028            :out std_logic;
     out2029            :out std_logic;
     out2030            :out std_logic;
     out2031            :out std_logic;
     out2032            :out std_logic;
     out2033            :out std_logic;
     out2034            :out std_logic;
     out2035            :out std_logic;
     out2036            :out std_logic;
     out2037            :out std_logic;
     out2038            :out std_logic;
     out2039            :out std_logic;
     out2040            :out std_logic;
     out2041            :out std_logic;
     out2042            :out std_logic;
     out2043            :out std_logic;
     out2044            :out std_logic;
     out2045            :out std_logic;
     out2046            :out std_logic;
     out2047            :out std_logic;
     out2048            :out std_logic;
     out2049            :out std_logic;
     out2050            :out std_logic;
     out2051            :out std_logic;
     out2052            :out std_logic;
     out2053            :out std_logic;
     out2054            :out std_logic;
     out2055            :out std_logic;
     out2056            :out std_logic;
     out2057            :out std_logic;
     out2058            :out std_logic;
     out2059            :out std_logic;
     out2060            :out std_logic;
     out2061            :out std_logic;
     out2062            :out std_logic;
     out2063            :out std_logic;
     out2064            :out std_logic;
     out2065            :out std_logic;
     out2066            :out std_logic;
     out2067            :out std_logic;
     out2068            :out std_logic;
     out2069            :out std_logic;
     out2070            :out std_logic;
     out2071            :out std_logic;
     out2072            :out std_logic;
     out2073            :out std_logic;
     out2074            :out std_logic;
     out2075            :out std_logic;
     out2076            :out std_logic;
     out2077            :out std_logic;
     out2078            :out std_logic;
     out2079            :out std_logic;
     out2080            :out std_logic;
     out2081            :out std_logic;
     out2082            :out std_logic;
     out2083            :out std_logic;
     out2084            :out std_logic;
     out2085            :out std_logic;
     out2086            :out std_logic;
     out2087            :out std_logic;
     out2088            :out std_logic;
     out2089            :out std_logic;
     out2090            :out std_logic;
     out2091            :out std_logic;
     out2092            :out std_logic;
     out2093            :out std_logic;
     out2094            :out std_logic;
     out2095            :out std_logic;
     out2096            :out std_logic;
     out2097            :out std_logic;
     out2098            :out std_logic;
     out2099            :out std_logic;
     out2100            :out std_logic;
     out2101            :out std_logic;
     out2102            :out std_logic;
     out2103            :out std_logic;
     out2104            :out std_logic;
     out2105            :out std_logic;
     out2106            :out std_logic;
     out2107            :out std_logic;
     out2108            :out std_logic;
     out2109            :out std_logic;
     out2110            :out std_logic;
     out2111            :out std_logic;
     out2112            :out std_logic;
     out2113            :out std_logic;
     out2114            :out std_logic;
     out2115            :out std_logic;
     out2116            :out std_logic;
     out2117            :out std_logic;
     out2118            :out std_logic;
     out2119            :out std_logic;
     out2120            :out std_logic;
     out2121            :out std_logic;
     out2122            :out std_logic;
     out2123            :out std_logic;
     out2124            :out std_logic;
     out2125            :out std_logic;
     out2126            :out std_logic;
     out2127            :out std_logic;
     out2128            :out std_logic;
     out2129            :out std_logic;
     out2130            :out std_logic;
     out2131            :out std_logic;
     out2132            :out std_logic;
     out2133            :out std_logic;
     out2134            :out std_logic;
     out2135            :out std_logic;
     out2136            :out std_logic;
     out2137            :out std_logic;
     out2138            :out std_logic;
     out2139            :out std_logic;
     out2140            :out std_logic;
     out2141            :out std_logic;
     out2142            :out std_logic;
     out2143            :out std_logic;
     out2144            :out std_logic;
     out2145            :out std_logic;
     out2146            :out std_logic;
     out2147            :out std_logic;
     out2148            :out std_logic;
     out2149            :out std_logic;
     out2150            :out std_logic;
     out2151            :out std_logic;
     out2152            :out std_logic;
     out2153            :out std_logic;
     out2154            :out std_logic;
     out2155            :out std_logic;
     out2156            :out std_logic;
     out2157            :out std_logic;
     out2158            :out std_logic;
     out2159            :out std_logic;
     out2160            :out std_logic;
     out2161            :out std_logic;
     out2162            :out std_logic;
     out2163            :out std_logic;
     out2164            :out std_logic;
     out2165            :out std_logic;
     out2166            :out std_logic;
     out2167            :out std_logic;
     out2168            :out std_logic;
     out2169            :out std_logic;
     out2170            :out std_logic;
     out2171            :out std_logic;
     out2172            :out std_logic;
     out2173            :out std_logic;
     out2174            :out std_logic;
     out2175            :out std_logic;
     out2176            :out std_logic;
     out2177            :out std_logic;
     out2178            :out std_logic;
     out2179            :out std_logic;
     out2180            :out std_logic;
     out2181            :out std_logic;
     out2182            :out std_logic;
     out2183            :out std_logic;
     out2184            :out std_logic;
     out2185            :out std_logic;
     out2186            :out std_logic;
     out2187            :out std_logic;
     out2188            :out std_logic;
     out2189            :out std_logic;
     out2190            :out std_logic;
     out2191            :out std_logic;
     out2192            :out std_logic;
     out2193            :out std_logic;
     out2194            :out std_logic;
     out2195            :out std_logic;
     out2196            :out std_logic;
     out2197            :out std_logic;
     out2198            :out std_logic;
     out2199            :out std_logic;
     out2200            :out std_logic;
     out2201            :out std_logic;
     out2202            :out std_logic;
     out2203            :out std_logic;
     out2204            :out std_logic;
     out2205            :out std_logic;
     out2206            :out std_logic;
     out2207            :out std_logic;
     out2208            :out std_logic;
     out2209            :out std_logic;
     out2210            :out std_logic;
     out2211            :out std_logic;
     out2212            :out std_logic;
     out2213            :out std_logic;
     out2214            :out std_logic;
     out2215            :out std_logic;
     out2216            :out std_logic;
     out2217            :out std_logic;
     out2218            :out std_logic;
     out2219            :out std_logic;
     out2220            :out std_logic;
     out2221            :out std_logic;
     out2222            :out std_logic;
     out2223            :out std_logic;
     out2224            :out std_logic;
     out2225            :out std_logic;
     out2226            :out std_logic;
     out2227            :out std_logic;
     out2228            :out std_logic;
     out2229            :out std_logic;
     out2230            :out std_logic;
     out2231            :out std_logic;
     out2232            :out std_logic;
     out2233            :out std_logic;
     out2234            :out std_logic;
     out2235            :out std_logic;
     out2236            :out std_logic;
     out2237            :out std_logic;
     out2238            :out std_logic;
     out2239            :out std_logic;
     out2240            :out std_logic;
     out2241            :out std_logic;
     out2242            :out std_logic;
     out2243            :out std_logic;
     out2244            :out std_logic;
     out2245            :out std_logic;
     out2246            :out std_logic;
     out2247            :out std_logic;
     out2248            :out std_logic;
     out2249            :out std_logic;
     out2250            :out std_logic;
     out2251            :out std_logic;
     out2252            :out std_logic;
     out2253            :out std_logic;
     out2254            :out std_logic;
     out2255            :out std_logic;
     out2256            :out std_logic;
     out2257            :out std_logic;
     out2258            :out std_logic;
     out2259            :out std_logic;
     out2260            :out std_logic;
     out2261            :out std_logic;
     out2262            :out std_logic;
     out2263            :out std_logic;
     out2264            :out std_logic;
     out2265            :out std_logic;
     out2266            :out std_logic;
     out2267            :out std_logic;
     out2268            :out std_logic;
     out2269            :out std_logic;
     out2270            :out std_logic;
     out2271            :out std_logic;
     out2272            :out std_logic;
     out2273            :out std_logic;
     out2274            :out std_logic;
     out2275            :out std_logic;
     out2276            :out std_logic;
     out2277            :out std_logic;
     out2278            :out std_logic;
     out2279            :out std_logic;
     out2280            :out std_logic;
     out2281            :out std_logic;
     out2282            :out std_logic;
     out2283            :out std_logic;
     out2284            :out std_logic;
     out2285            :out std_logic;
     out2286            :out std_logic;
     out2287            :out std_logic;
     out2288            :out std_logic;
     out2289            :out std_logic;
     out2290            :out std_logic;
     out2291            :out std_logic;
     out2292            :out std_logic;
     out2293            :out std_logic;
     out2294            :out std_logic;
     out2295            :out std_logic;
     out2296            :out std_logic;
     out2297            :out std_logic;
     out2298            :out std_logic;
     out2299            :out std_logic;
     out2300            :out std_logic;
     out2301            :out std_logic;
     out2302            :out std_logic;
     out2303            :out std_logic;
     out2304            :out std_logic;
     end_cnt,end_vnt      :out std_logic
);
END;
ARCHITECTURE ldpc_arch OF ldpc IS
------------------------VNPU3_3 Component--------------------------------------
COMPONENT VNPU3_3 is PORT(
start_vn_3                        :   IN    std_logic;
clk                               :   IN    std_logic;
rst                               :   IN    std_logic;
Lc_3                              :   IN    std_logic_vector(8 DOWNTO 0);
L1_3                              :   IN    std_logic_vector(8 DOWNTO 0);
L2_3                              :   IN    std_logic_vector(8 DOWNTO 0);
L3_3                              :   IN    std_logic_vector(8 DOWNTO 0);
Z1_3                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z2_3                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z3_3                              :   OUT    std_logic_vector(8 DOWNTO 0);
SI_3                              :   OUT    std_logic;
end_vn_3                          :   OUT    std_logic);
 end component;
------------------------VNPU6_6 Component--------------------------------------
COMPONENT VNPU6_6 is PORT(
start_vn_6                        :   IN    std_logic;
clk                               :   IN    std_logic;
rst                               :   IN    std_logic;
Lc_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L1_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L2_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L3_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L4_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L5_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L6_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z1_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z2_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z3_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z4_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z5_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z6_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
SI_6                              :   OUT    std_logic;
end_vn_6                          :   OUT    std_logic);
 end component;
------------------------VNPU2_2 Component--------------------------------------
COMPONENT VNPU2_2 is PORT(
start_vn_2                        :   IN    std_logic;
clk                               :   IN    std_logic;
rst                               :   IN    std_logic;
Lc_2                              :   IN    std_logic_vector(8 DOWNTO 0);
L1_2                              :   IN    std_logic_vector(8 DOWNTO 0);
L2_2                              :   IN    std_logic_vector(8 DOWNTO 0);
Z1_2                              :   OUT    std_logic_vector(8 DOWNTO 0);
Z2_2                              :   OUT    std_logic_vector(8 DOWNTO 0);
SI_2                              :   OUT    std_logic;
end_vn_2                          :   OUT    std_logic);
 end component;
---------------------CNPU6_6 Component---------------------------------------------------
COMPONENT CNPU6_6 is PORT(
start_cn_6                        :   IN    std_logic;
clk                               :   IN    std_logic;
rst                               :   IN    std_logic;
Z1_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z2_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z3_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z4_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z5_6                              :   IN    std_logic_vector(8 DOWNTO 0);
Z6_6                              :   IN    std_logic_vector(8 DOWNTO 0);
L1_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
L2_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
L3_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
L4_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
L5_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
L6_6                              :   OUT    std_logic_vector(8 DOWNTO 0);
end_cn_6                          :   OUT    std_logic);
 end component;
---------------------CNPU7_7 Component---------------------------------------------------
COMPONENT CNPU7_7 is PORT(
start_cn_7                        :   IN    std_logic;
clk                               :   IN    std_logic;
rst                               :   IN    std_logic;
Z1_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z2_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z3_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z4_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z5_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z6_7                              :   IN    std_logic_vector(8 DOWNTO 0);
Z7_7                              :   IN    std_logic_vector(8 DOWNTO 0);
L1_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L2_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L3_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L4_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L5_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L6_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
L7_7                              :   OUT    std_logic_vector(8 DOWNTO 0);
end_cn_7                          :   OUT    std_logic);
 end component;
FOR ALL : VNPU3_3
USE ENTITY work.VNPU3_3(rtl);
FOR ALL : VNPU6_6
USE ENTITY work.VNPU6_6(rtl);
FOR ALL : VNPU2_2
USE ENTITY work.VNPU2_2(rtl);
FOR ALL : CNPU6_6
USE ENTITY work.CNPU6_6(rtl);
FOR ALL : CNPU7_7
USE ENTITY work.CNPU7_7(rtl);
signal V191C1,V266C1,V824C1,V948C1,V1160C1,V1249C1,C1V191,C1V266,C1V824,C1V948,C1V1160,C1V1249:std_logic_vector(8 downto 0);
signal V192C2,V267C2,V825C2,V949C2,V1161C2,V1250C2,C2V192,C2V267,C2V825,C2V949,C2V1161,C2V1250:std_logic_vector(8 downto 0);
signal V97C3,V268C3,V826C3,V950C3,V1162C3,V1251C3,C3V97,C3V268,C3V826,C3V950,C3V1162,C3V1251:std_logic_vector(8 downto 0);
signal V98C4,V269C4,V827C4,V951C4,V1163C4,V1252C4,C4V98,C4V269,C4V827,C4V951,C4V1163,C4V1252:std_logic_vector(8 downto 0);
signal V99C5,V270C5,V828C5,V952C5,V1164C5,V1253C5,C5V99,C5V270,C5V828,C5V952,C5V1164,C5V1253:std_logic_vector(8 downto 0);
signal V100C6,V271C6,V829C6,V953C6,V1165C6,V1254C6,C6V100,C6V271,C6V829,C6V953,C6V1165,C6V1254:std_logic_vector(8 downto 0);
signal V101C7,V272C7,V830C7,V954C7,V1166C7,V1255C7,C7V101,C7V272,C7V830,C7V954,C7V1166,C7V1255:std_logic_vector(8 downto 0);
signal V102C8,V273C8,V831C8,V955C8,V1167C8,V1256C8,C8V102,C8V273,C8V831,C8V955,C8V1167,C8V1256:std_logic_vector(8 downto 0);
signal V103C9,V274C9,V832C9,V956C9,V1168C9,V1257C9,C9V103,C9V274,C9V832,C9V956,C9V1168,C9V1257:std_logic_vector(8 downto 0);
signal V104C10,V275C10,V833C10,V957C10,V1169C10,V1258C10,C10V104,C10V275,C10V833,C10V957,C10V1169,C10V1258:std_logic_vector(8 downto 0);
signal V105C11,V276C11,V834C11,V958C11,V1170C11,V1259C11,C11V105,C11V276,C11V834,C11V958,C11V1170,C11V1259:std_logic_vector(8 downto 0);
signal V106C12,V277C12,V835C12,V959C12,V1171C12,V1260C12,C12V106,C12V277,C12V835,C12V959,C12V1171,C12V1260:std_logic_vector(8 downto 0);
signal V107C13,V278C13,V836C13,V960C13,V1172C13,V1261C13,C13V107,C13V278,C13V836,C13V960,C13V1172,C13V1261:std_logic_vector(8 downto 0);
signal V108C14,V279C14,V837C14,V865C14,V1173C14,V1262C14,C14V108,C14V279,C14V837,C14V865,C14V1173,C14V1262:std_logic_vector(8 downto 0);
signal V109C15,V280C15,V838C15,V866C15,V1174C15,V1263C15,C15V109,C15V280,C15V838,C15V866,C15V1174,C15V1263:std_logic_vector(8 downto 0);
signal V110C16,V281C16,V839C16,V867C16,V1175C16,V1264C16,C16V110,C16V281,C16V839,C16V867,C16V1175,C16V1264:std_logic_vector(8 downto 0);
signal V111C17,V282C17,V840C17,V868C17,V1176C17,V1265C17,C17V111,C17V282,C17V840,C17V868,C17V1176,C17V1265:std_logic_vector(8 downto 0);
signal V112C18,V283C18,V841C18,V869C18,V1177C18,V1266C18,C18V112,C18V283,C18V841,C18V869,C18V1177,C18V1266:std_logic_vector(8 downto 0);
signal V113C19,V284C19,V842C19,V870C19,V1178C19,V1267C19,C19V113,C19V284,C19V842,C19V870,C19V1178,C19V1267:std_logic_vector(8 downto 0);
signal V114C20,V285C20,V843C20,V871C20,V1179C20,V1268C20,C20V114,C20V285,C20V843,C20V871,C20V1179,C20V1268:std_logic_vector(8 downto 0);
signal V115C21,V286C21,V844C21,V872C21,V1180C21,V1269C21,C21V115,C21V286,C21V844,C21V872,C21V1180,C21V1269:std_logic_vector(8 downto 0);
signal V116C22,V287C22,V845C22,V873C22,V1181C22,V1270C22,C22V116,C22V287,C22V845,C22V873,C22V1181,C22V1270:std_logic_vector(8 downto 0);
signal V117C23,V288C23,V846C23,V874C23,V1182C23,V1271C23,C23V117,C23V288,C23V846,C23V874,C23V1182,C23V1271:std_logic_vector(8 downto 0);
signal V118C24,V193C24,V847C24,V875C24,V1183C24,V1272C24,C24V118,C24V193,C24V847,C24V875,C24V1183,C24V1272:std_logic_vector(8 downto 0);
signal V119C25,V194C25,V848C25,V876C25,V1184C25,V1273C25,C25V119,C25V194,C25V848,C25V876,C25V1184,C25V1273:std_logic_vector(8 downto 0);
signal V120C26,V195C26,V849C26,V877C26,V1185C26,V1274C26,C26V120,C26V195,C26V849,C26V877,C26V1185,C26V1274:std_logic_vector(8 downto 0);
signal V121C27,V196C27,V850C27,V878C27,V1186C27,V1275C27,C27V121,C27V196,C27V850,C27V878,C27V1186,C27V1275:std_logic_vector(8 downto 0);
signal V122C28,V197C28,V851C28,V879C28,V1187C28,V1276C28,C28V122,C28V197,C28V851,C28V879,C28V1187,C28V1276:std_logic_vector(8 downto 0);
signal V123C29,V198C29,V852C29,V880C29,V1188C29,V1277C29,C29V123,C29V198,C29V852,C29V880,C29V1188,C29V1277:std_logic_vector(8 downto 0);
signal V124C30,V199C30,V853C30,V881C30,V1189C30,V1278C30,C30V124,C30V199,C30V853,C30V881,C30V1189,C30V1278:std_logic_vector(8 downto 0);
signal V125C31,V200C31,V854C31,V882C31,V1190C31,V1279C31,C31V125,C31V200,C31V854,C31V882,C31V1190,C31V1279:std_logic_vector(8 downto 0);
signal V126C32,V201C32,V855C32,V883C32,V1191C32,V1280C32,C32V126,C32V201,C32V855,C32V883,C32V1191,C32V1280:std_logic_vector(8 downto 0);
signal V127C33,V202C33,V856C33,V884C33,V1192C33,V1281C33,C33V127,C33V202,C33V856,C33V884,C33V1192,C33V1281:std_logic_vector(8 downto 0);
signal V128C34,V203C34,V857C34,V885C34,V1193C34,V1282C34,C34V128,C34V203,C34V857,C34V885,C34V1193,C34V1282:std_logic_vector(8 downto 0);
signal V129C35,V204C35,V858C35,V886C35,V1194C35,V1283C35,C35V129,C35V204,C35V858,C35V886,C35V1194,C35V1283:std_logic_vector(8 downto 0);
signal V130C36,V205C36,V859C36,V887C36,V1195C36,V1284C36,C36V130,C36V205,C36V859,C36V887,C36V1195,C36V1284:std_logic_vector(8 downto 0);
signal V131C37,V206C37,V860C37,V888C37,V1196C37,V1285C37,C37V131,C37V206,C37V860,C37V888,C37V1196,C37V1285:std_logic_vector(8 downto 0);
signal V132C38,V207C38,V861C38,V889C38,V1197C38,V1286C38,C38V132,C38V207,C38V861,C38V889,C38V1197,C38V1286:std_logic_vector(8 downto 0);
signal V133C39,V208C39,V862C39,V890C39,V1198C39,V1287C39,C39V133,C39V208,C39V862,C39V890,C39V1198,C39V1287:std_logic_vector(8 downto 0);
signal V134C40,V209C40,V863C40,V891C40,V1199C40,V1288C40,C40V134,C40V209,C40V863,C40V891,C40V1199,C40V1288:std_logic_vector(8 downto 0);
signal V135C41,V210C41,V864C41,V892C41,V1200C41,V1289C41,C41V135,C41V210,C41V864,C41V892,C41V1200,C41V1289:std_logic_vector(8 downto 0);
signal V136C42,V211C42,V769C42,V893C42,V1201C42,V1290C42,C42V136,C42V211,C42V769,C42V893,C42V1201,C42V1290:std_logic_vector(8 downto 0);
signal V137C43,V212C43,V770C43,V894C43,V1202C43,V1291C43,C43V137,C43V212,C43V770,C43V894,C43V1202,C43V1291:std_logic_vector(8 downto 0);
signal V138C44,V213C44,V771C44,V895C44,V1203C44,V1292C44,C44V138,C44V213,C44V771,C44V895,C44V1203,C44V1292:std_logic_vector(8 downto 0);
signal V139C45,V214C45,V772C45,V896C45,V1204C45,V1293C45,C45V139,C45V214,C45V772,C45V896,C45V1204,C45V1293:std_logic_vector(8 downto 0);
signal V140C46,V215C46,V773C46,V897C46,V1205C46,V1294C46,C46V140,C46V215,C46V773,C46V897,C46V1205,C46V1294:std_logic_vector(8 downto 0);
signal V141C47,V216C47,V774C47,V898C47,V1206C47,V1295C47,C47V141,C47V216,C47V774,C47V898,C47V1206,C47V1295:std_logic_vector(8 downto 0);
signal V142C48,V217C48,V775C48,V899C48,V1207C48,V1296C48,C48V142,C48V217,C48V775,C48V899,C48V1207,C48V1296:std_logic_vector(8 downto 0);
signal V143C49,V218C49,V776C49,V900C49,V1208C49,V1297C49,C49V143,C49V218,C49V776,C49V900,C49V1208,C49V1297:std_logic_vector(8 downto 0);
signal V144C50,V219C50,V777C50,V901C50,V1209C50,V1298C50,C50V144,C50V219,C50V777,C50V901,C50V1209,C50V1298:std_logic_vector(8 downto 0);
signal V145C51,V220C51,V778C51,V902C51,V1210C51,V1299C51,C51V145,C51V220,C51V778,C51V902,C51V1210,C51V1299:std_logic_vector(8 downto 0);
signal V146C52,V221C52,V779C52,V903C52,V1211C52,V1300C52,C52V146,C52V221,C52V779,C52V903,C52V1211,C52V1300:std_logic_vector(8 downto 0);
signal V147C53,V222C53,V780C53,V904C53,V1212C53,V1301C53,C53V147,C53V222,C53V780,C53V904,C53V1212,C53V1301:std_logic_vector(8 downto 0);
signal V148C54,V223C54,V781C54,V905C54,V1213C54,V1302C54,C54V148,C54V223,C54V781,C54V905,C54V1213,C54V1302:std_logic_vector(8 downto 0);
signal V149C55,V224C55,V782C55,V906C55,V1214C55,V1303C55,C55V149,C55V224,C55V782,C55V906,C55V1214,C55V1303:std_logic_vector(8 downto 0);
signal V150C56,V225C56,V783C56,V907C56,V1215C56,V1304C56,C56V150,C56V225,C56V783,C56V907,C56V1215,C56V1304:std_logic_vector(8 downto 0);
signal V151C57,V226C57,V784C57,V908C57,V1216C57,V1305C57,C57V151,C57V226,C57V784,C57V908,C57V1216,C57V1305:std_logic_vector(8 downto 0);
signal V152C58,V227C58,V785C58,V909C58,V1217C58,V1306C58,C58V152,C58V227,C58V785,C58V909,C58V1217,C58V1306:std_logic_vector(8 downto 0);
signal V153C59,V228C59,V786C59,V910C59,V1218C59,V1307C59,C59V153,C59V228,C59V786,C59V910,C59V1218,C59V1307:std_logic_vector(8 downto 0);
signal V154C60,V229C60,V787C60,V911C60,V1219C60,V1308C60,C60V154,C60V229,C60V787,C60V911,C60V1219,C60V1308:std_logic_vector(8 downto 0);
signal V155C61,V230C61,V788C61,V912C61,V1220C61,V1309C61,C61V155,C61V230,C61V788,C61V912,C61V1220,C61V1309:std_logic_vector(8 downto 0);
signal V156C62,V231C62,V789C62,V913C62,V1221C62,V1310C62,C62V156,C62V231,C62V789,C62V913,C62V1221,C62V1310:std_logic_vector(8 downto 0);
signal V157C63,V232C63,V790C63,V914C63,V1222C63,V1311C63,C63V157,C63V232,C63V790,C63V914,C63V1222,C63V1311:std_logic_vector(8 downto 0);
signal V158C64,V233C64,V791C64,V915C64,V1223C64,V1312C64,C64V158,C64V233,C64V791,C64V915,C64V1223,C64V1312:std_logic_vector(8 downto 0);
signal V159C65,V234C65,V792C65,V916C65,V1224C65,V1313C65,C65V159,C65V234,C65V792,C65V916,C65V1224,C65V1313:std_logic_vector(8 downto 0);
signal V160C66,V235C66,V793C66,V917C66,V1225C66,V1314C66,C66V160,C66V235,C66V793,C66V917,C66V1225,C66V1314:std_logic_vector(8 downto 0);
signal V161C67,V236C67,V794C67,V918C67,V1226C67,V1315C67,C67V161,C67V236,C67V794,C67V918,C67V1226,C67V1315:std_logic_vector(8 downto 0);
signal V162C68,V237C68,V795C68,V919C68,V1227C68,V1316C68,C68V162,C68V237,C68V795,C68V919,C68V1227,C68V1316:std_logic_vector(8 downto 0);
signal V163C69,V238C69,V796C69,V920C69,V1228C69,V1317C69,C69V163,C69V238,C69V796,C69V920,C69V1228,C69V1317:std_logic_vector(8 downto 0);
signal V164C70,V239C70,V797C70,V921C70,V1229C70,V1318C70,C70V164,C70V239,C70V797,C70V921,C70V1229,C70V1318:std_logic_vector(8 downto 0);
signal V165C71,V240C71,V798C71,V922C71,V1230C71,V1319C71,C71V165,C71V240,C71V798,C71V922,C71V1230,C71V1319:std_logic_vector(8 downto 0);
signal V166C72,V241C72,V799C72,V923C72,V1231C72,V1320C72,C72V166,C72V241,C72V799,C72V923,C72V1231,C72V1320:std_logic_vector(8 downto 0);
signal V167C73,V242C73,V800C73,V924C73,V1232C73,V1321C73,C73V167,C73V242,C73V800,C73V924,C73V1232,C73V1321:std_logic_vector(8 downto 0);
signal V168C74,V243C74,V801C74,V925C74,V1233C74,V1322C74,C74V168,C74V243,C74V801,C74V925,C74V1233,C74V1322:std_logic_vector(8 downto 0);
signal V169C75,V244C75,V802C75,V926C75,V1234C75,V1323C75,C75V169,C75V244,C75V802,C75V926,C75V1234,C75V1323:std_logic_vector(8 downto 0);
signal V170C76,V245C76,V803C76,V927C76,V1235C76,V1324C76,C76V170,C76V245,C76V803,C76V927,C76V1235,C76V1324:std_logic_vector(8 downto 0);
signal V171C77,V246C77,V804C77,V928C77,V1236C77,V1325C77,C77V171,C77V246,C77V804,C77V928,C77V1236,C77V1325:std_logic_vector(8 downto 0);
signal V172C78,V247C78,V805C78,V929C78,V1237C78,V1326C78,C78V172,C78V247,C78V805,C78V929,C78V1237,C78V1326:std_logic_vector(8 downto 0);
signal V173C79,V248C79,V806C79,V930C79,V1238C79,V1327C79,C79V173,C79V248,C79V806,C79V930,C79V1238,C79V1327:std_logic_vector(8 downto 0);
signal V174C80,V249C80,V807C80,V931C80,V1239C80,V1328C80,C80V174,C80V249,C80V807,C80V931,C80V1239,C80V1328:std_logic_vector(8 downto 0);
signal V175C81,V250C81,V808C81,V932C81,V1240C81,V1329C81,C81V175,C81V250,C81V808,C81V932,C81V1240,C81V1329:std_logic_vector(8 downto 0);
signal V176C82,V251C82,V809C82,V933C82,V1241C82,V1330C82,C82V176,C82V251,C82V809,C82V933,C82V1241,C82V1330:std_logic_vector(8 downto 0);
signal V177C83,V252C83,V810C83,V934C83,V1242C83,V1331C83,C83V177,C83V252,C83V810,C83V934,C83V1242,C83V1331:std_logic_vector(8 downto 0);
signal V178C84,V253C84,V811C84,V935C84,V1243C84,V1332C84,C84V178,C84V253,C84V811,C84V935,C84V1243,C84V1332:std_logic_vector(8 downto 0);
signal V179C85,V254C85,V812C85,V936C85,V1244C85,V1333C85,C85V179,C85V254,C85V812,C85V936,C85V1244,C85V1333:std_logic_vector(8 downto 0);
signal V180C86,V255C86,V813C86,V937C86,V1245C86,V1334C86,C86V180,C86V255,C86V813,C86V937,C86V1245,C86V1334:std_logic_vector(8 downto 0);
signal V181C87,V256C87,V814C87,V938C87,V1246C87,V1335C87,C87V181,C87V256,C87V814,C87V938,C87V1246,C87V1335:std_logic_vector(8 downto 0);
signal V182C88,V257C88,V815C88,V939C88,V1247C88,V1336C88,C88V182,C88V257,C88V815,C88V939,C88V1247,C88V1336:std_logic_vector(8 downto 0);
signal V183C89,V258C89,V816C89,V940C89,V1248C89,V1337C89,C89V183,C89V258,C89V816,C89V940,C89V1248,C89V1337:std_logic_vector(8 downto 0);
signal V184C90,V259C90,V817C90,V941C90,V1153C90,V1338C90,C90V184,C90V259,C90V817,C90V941,C90V1153,C90V1338:std_logic_vector(8 downto 0);
signal V185C91,V260C91,V818C91,V942C91,V1154C91,V1339C91,C91V185,C91V260,C91V818,C91V942,C91V1154,C91V1339:std_logic_vector(8 downto 0);
signal V186C92,V261C92,V819C92,V943C92,V1155C92,V1340C92,C92V186,C92V261,C92V819,C92V943,C92V1155,C92V1340:std_logic_vector(8 downto 0);
signal V187C93,V262C93,V820C93,V944C93,V1156C93,V1341C93,C93V187,C93V262,C93V820,C93V944,C93V1156,C93V1341:std_logic_vector(8 downto 0);
signal V188C94,V263C94,V821C94,V945C94,V1157C94,V1342C94,C94V188,C94V263,C94V821,C94V945,C94V1157,C94V1342:std_logic_vector(8 downto 0);
signal V189C95,V264C95,V822C95,V946C95,V1158C95,V1343C95,C95V189,C95V264,C95V822,C95V946,C95V1158,C95V1343:std_logic_vector(8 downto 0);
signal V190C96,V265C96,V823C96,V947C96,V1159C96,V1344C96,C96V190,C96V265,C96V823,C96V947,C96V1159,C96V1344:std_logic_vector(8 downto 0);
signal V124C97,V503C97,V656C97,V682C97,V1069C97,V1249C97,V1345C97,C97V124,C97V503,C97V656,C97V682,C97V1069,C97V1249,C97V1345:std_logic_vector(8 downto 0);
signal V125C98,V504C98,V657C98,V683C98,V1070C98,V1250C98,V1346C98,C98V125,C98V504,C98V657,C98V683,C98V1070,C98V1250,C98V1346:std_logic_vector(8 downto 0);
signal V126C99,V505C99,V658C99,V684C99,V1071C99,V1251C99,V1347C99,C99V126,C99V505,C99V658,C99V684,C99V1071,C99V1251,C99V1347:std_logic_vector(8 downto 0);
signal V127C100,V506C100,V659C100,V685C100,V1072C100,V1252C100,V1348C100,C100V127,C100V506,C100V659,C100V685,C100V1072,C100V1252,C100V1348:std_logic_vector(8 downto 0);
signal V128C101,V507C101,V660C101,V686C101,V1073C101,V1253C101,V1349C101,C101V128,C101V507,C101V660,C101V686,C101V1073,C101V1253,C101V1349:std_logic_vector(8 downto 0);
signal V129C102,V508C102,V661C102,V687C102,V1074C102,V1254C102,V1350C102,C102V129,C102V508,C102V661,C102V687,C102V1074,C102V1254,C102V1350:std_logic_vector(8 downto 0);
signal V130C103,V509C103,V662C103,V688C103,V1075C103,V1255C103,V1351C103,C103V130,C103V509,C103V662,C103V688,C103V1075,C103V1255,C103V1351:std_logic_vector(8 downto 0);
signal V131C104,V510C104,V663C104,V689C104,V1076C104,V1256C104,V1352C104,C104V131,C104V510,C104V663,C104V689,C104V1076,C104V1256,C104V1352:std_logic_vector(8 downto 0);
signal V132C105,V511C105,V664C105,V690C105,V1077C105,V1257C105,V1353C105,C105V132,C105V511,C105V664,C105V690,C105V1077,C105V1257,C105V1353:std_logic_vector(8 downto 0);
signal V133C106,V512C106,V665C106,V691C106,V1078C106,V1258C106,V1354C106,C106V133,C106V512,C106V665,C106V691,C106V1078,C106V1258,C106V1354:std_logic_vector(8 downto 0);
signal V134C107,V513C107,V666C107,V692C107,V1079C107,V1259C107,V1355C107,C107V134,C107V513,C107V666,C107V692,C107V1079,C107V1259,C107V1355:std_logic_vector(8 downto 0);
signal V135C108,V514C108,V667C108,V693C108,V1080C108,V1260C108,V1356C108,C108V135,C108V514,C108V667,C108V693,C108V1080,C108V1260,C108V1356:std_logic_vector(8 downto 0);
signal V136C109,V515C109,V668C109,V694C109,V1081C109,V1261C109,V1357C109,C109V136,C109V515,C109V668,C109V694,C109V1081,C109V1261,C109V1357:std_logic_vector(8 downto 0);
signal V137C110,V516C110,V669C110,V695C110,V1082C110,V1262C110,V1358C110,C110V137,C110V516,C110V669,C110V695,C110V1082,C110V1262,C110V1358:std_logic_vector(8 downto 0);
signal V138C111,V517C111,V670C111,V696C111,V1083C111,V1263C111,V1359C111,C111V138,C111V517,C111V670,C111V696,C111V1083,C111V1263,C111V1359:std_logic_vector(8 downto 0);
signal V139C112,V518C112,V671C112,V697C112,V1084C112,V1264C112,V1360C112,C112V139,C112V518,C112V671,C112V697,C112V1084,C112V1264,C112V1360:std_logic_vector(8 downto 0);
signal V140C113,V519C113,V672C113,V698C113,V1085C113,V1265C113,V1361C113,C113V140,C113V519,C113V672,C113V698,C113V1085,C113V1265,C113V1361:std_logic_vector(8 downto 0);
signal V141C114,V520C114,V577C114,V699C114,V1086C114,V1266C114,V1362C114,C114V141,C114V520,C114V577,C114V699,C114V1086,C114V1266,C114V1362:std_logic_vector(8 downto 0);
signal V142C115,V521C115,V578C115,V700C115,V1087C115,V1267C115,V1363C115,C115V142,C115V521,C115V578,C115V700,C115V1087,C115V1267,C115V1363:std_logic_vector(8 downto 0);
signal V143C116,V522C116,V579C116,V701C116,V1088C116,V1268C116,V1364C116,C116V143,C116V522,C116V579,C116V701,C116V1088,C116V1268,C116V1364:std_logic_vector(8 downto 0);
signal V144C117,V523C117,V580C117,V702C117,V1089C117,V1269C117,V1365C117,C117V144,C117V523,C117V580,C117V702,C117V1089,C117V1269,C117V1365:std_logic_vector(8 downto 0);
signal V145C118,V524C118,V581C118,V703C118,V1090C118,V1270C118,V1366C118,C118V145,C118V524,C118V581,C118V703,C118V1090,C118V1270,C118V1366:std_logic_vector(8 downto 0);
signal V146C119,V525C119,V582C119,V704C119,V1091C119,V1271C119,V1367C119,C119V146,C119V525,C119V582,C119V704,C119V1091,C119V1271,C119V1367:std_logic_vector(8 downto 0);
signal V147C120,V526C120,V583C120,V705C120,V1092C120,V1272C120,V1368C120,C120V147,C120V526,C120V583,C120V705,C120V1092,C120V1272,C120V1368:std_logic_vector(8 downto 0);
signal V148C121,V527C121,V584C121,V706C121,V1093C121,V1273C121,V1369C121,C121V148,C121V527,C121V584,C121V706,C121V1093,C121V1273,C121V1369:std_logic_vector(8 downto 0);
signal V149C122,V528C122,V585C122,V707C122,V1094C122,V1274C122,V1370C122,C122V149,C122V528,C122V585,C122V707,C122V1094,C122V1274,C122V1370:std_logic_vector(8 downto 0);
signal V150C123,V529C123,V586C123,V708C123,V1095C123,V1275C123,V1371C123,C123V150,C123V529,C123V586,C123V708,C123V1095,C123V1275,C123V1371:std_logic_vector(8 downto 0);
signal V151C124,V530C124,V587C124,V709C124,V1096C124,V1276C124,V1372C124,C124V151,C124V530,C124V587,C124V709,C124V1096,C124V1276,C124V1372:std_logic_vector(8 downto 0);
signal V152C125,V531C125,V588C125,V710C125,V1097C125,V1277C125,V1373C125,C125V152,C125V531,C125V588,C125V710,C125V1097,C125V1277,C125V1373:std_logic_vector(8 downto 0);
signal V153C126,V532C126,V589C126,V711C126,V1098C126,V1278C126,V1374C126,C126V153,C126V532,C126V589,C126V711,C126V1098,C126V1278,C126V1374:std_logic_vector(8 downto 0);
signal V154C127,V533C127,V590C127,V712C127,V1099C127,V1279C127,V1375C127,C127V154,C127V533,C127V590,C127V712,C127V1099,C127V1279,C127V1375:std_logic_vector(8 downto 0);
signal V155C128,V534C128,V591C128,V713C128,V1100C128,V1280C128,V1376C128,C128V155,C128V534,C128V591,C128V713,C128V1100,C128V1280,C128V1376:std_logic_vector(8 downto 0);
signal V156C129,V535C129,V592C129,V714C129,V1101C129,V1281C129,V1377C129,C129V156,C129V535,C129V592,C129V714,C129V1101,C129V1281,C129V1377:std_logic_vector(8 downto 0);
signal V157C130,V536C130,V593C130,V715C130,V1102C130,V1282C130,V1378C130,C130V157,C130V536,C130V593,C130V715,C130V1102,C130V1282,C130V1378:std_logic_vector(8 downto 0);
signal V158C131,V537C131,V594C131,V716C131,V1103C131,V1283C131,V1379C131,C131V158,C131V537,C131V594,C131V716,C131V1103,C131V1283,C131V1379:std_logic_vector(8 downto 0);
signal V159C132,V538C132,V595C132,V717C132,V1104C132,V1284C132,V1380C132,C132V159,C132V538,C132V595,C132V717,C132V1104,C132V1284,C132V1380:std_logic_vector(8 downto 0);
signal V160C133,V539C133,V596C133,V718C133,V1105C133,V1285C133,V1381C133,C133V160,C133V539,C133V596,C133V718,C133V1105,C133V1285,C133V1381:std_logic_vector(8 downto 0);
signal V161C134,V540C134,V597C134,V719C134,V1106C134,V1286C134,V1382C134,C134V161,C134V540,C134V597,C134V719,C134V1106,C134V1286,C134V1382:std_logic_vector(8 downto 0);
signal V162C135,V541C135,V598C135,V720C135,V1107C135,V1287C135,V1383C135,C135V162,C135V541,C135V598,C135V720,C135V1107,C135V1287,C135V1383:std_logic_vector(8 downto 0);
signal V163C136,V542C136,V599C136,V721C136,V1108C136,V1288C136,V1384C136,C136V163,C136V542,C136V599,C136V721,C136V1108,C136V1288,C136V1384:std_logic_vector(8 downto 0);
signal V164C137,V543C137,V600C137,V722C137,V1109C137,V1289C137,V1385C137,C137V164,C137V543,C137V600,C137V722,C137V1109,C137V1289,C137V1385:std_logic_vector(8 downto 0);
signal V165C138,V544C138,V601C138,V723C138,V1110C138,V1290C138,V1386C138,C138V165,C138V544,C138V601,C138V723,C138V1110,C138V1290,C138V1386:std_logic_vector(8 downto 0);
signal V166C139,V545C139,V602C139,V724C139,V1111C139,V1291C139,V1387C139,C139V166,C139V545,C139V602,C139V724,C139V1111,C139V1291,C139V1387:std_logic_vector(8 downto 0);
signal V167C140,V546C140,V603C140,V725C140,V1112C140,V1292C140,V1388C140,C140V167,C140V546,C140V603,C140V725,C140V1112,C140V1292,C140V1388:std_logic_vector(8 downto 0);
signal V168C141,V547C141,V604C141,V726C141,V1113C141,V1293C141,V1389C141,C141V168,C141V547,C141V604,C141V726,C141V1113,C141V1293,C141V1389:std_logic_vector(8 downto 0);
signal V169C142,V548C142,V605C142,V727C142,V1114C142,V1294C142,V1390C142,C142V169,C142V548,C142V605,C142V727,C142V1114,C142V1294,C142V1390:std_logic_vector(8 downto 0);
signal V170C143,V549C143,V606C143,V728C143,V1115C143,V1295C143,V1391C143,C143V170,C143V549,C143V606,C143V728,C143V1115,C143V1295,C143V1391:std_logic_vector(8 downto 0);
signal V171C144,V550C144,V607C144,V729C144,V1116C144,V1296C144,V1392C144,C144V171,C144V550,C144V607,C144V729,C144V1116,C144V1296,C144V1392:std_logic_vector(8 downto 0);
signal V172C145,V551C145,V608C145,V730C145,V1117C145,V1297C145,V1393C145,C145V172,C145V551,C145V608,C145V730,C145V1117,C145V1297,C145V1393:std_logic_vector(8 downto 0);
signal V173C146,V552C146,V609C146,V731C146,V1118C146,V1298C146,V1394C146,C146V173,C146V552,C146V609,C146V731,C146V1118,C146V1298,C146V1394:std_logic_vector(8 downto 0);
signal V174C147,V553C147,V610C147,V732C147,V1119C147,V1299C147,V1395C147,C147V174,C147V553,C147V610,C147V732,C147V1119,C147V1299,C147V1395:std_logic_vector(8 downto 0);
signal V175C148,V554C148,V611C148,V733C148,V1120C148,V1300C148,V1396C148,C148V175,C148V554,C148V611,C148V733,C148V1120,C148V1300,C148V1396:std_logic_vector(8 downto 0);
signal V176C149,V555C149,V612C149,V734C149,V1121C149,V1301C149,V1397C149,C149V176,C149V555,C149V612,C149V734,C149V1121,C149V1301,C149V1397:std_logic_vector(8 downto 0);
signal V177C150,V556C150,V613C150,V735C150,V1122C150,V1302C150,V1398C150,C150V177,C150V556,C150V613,C150V735,C150V1122,C150V1302,C150V1398:std_logic_vector(8 downto 0);
signal V178C151,V557C151,V614C151,V736C151,V1123C151,V1303C151,V1399C151,C151V178,C151V557,C151V614,C151V736,C151V1123,C151V1303,C151V1399:std_logic_vector(8 downto 0);
signal V179C152,V558C152,V615C152,V737C152,V1124C152,V1304C152,V1400C152,C152V179,C152V558,C152V615,C152V737,C152V1124,C152V1304,C152V1400:std_logic_vector(8 downto 0);
signal V180C153,V559C153,V616C153,V738C153,V1125C153,V1305C153,V1401C153,C153V180,C153V559,C153V616,C153V738,C153V1125,C153V1305,C153V1401:std_logic_vector(8 downto 0);
signal V181C154,V560C154,V617C154,V739C154,V1126C154,V1306C154,V1402C154,C154V181,C154V560,C154V617,C154V739,C154V1126,C154V1306,C154V1402:std_logic_vector(8 downto 0);
signal V182C155,V561C155,V618C155,V740C155,V1127C155,V1307C155,V1403C155,C155V182,C155V561,C155V618,C155V740,C155V1127,C155V1307,C155V1403:std_logic_vector(8 downto 0);
signal V183C156,V562C156,V619C156,V741C156,V1128C156,V1308C156,V1404C156,C156V183,C156V562,C156V619,C156V741,C156V1128,C156V1308,C156V1404:std_logic_vector(8 downto 0);
signal V184C157,V563C157,V620C157,V742C157,V1129C157,V1309C157,V1405C157,C157V184,C157V563,C157V620,C157V742,C157V1129,C157V1309,C157V1405:std_logic_vector(8 downto 0);
signal V185C158,V564C158,V621C158,V743C158,V1130C158,V1310C158,V1406C158,C158V185,C158V564,C158V621,C158V743,C158V1130,C158V1310,C158V1406:std_logic_vector(8 downto 0);
signal V186C159,V565C159,V622C159,V744C159,V1131C159,V1311C159,V1407C159,C159V186,C159V565,C159V622,C159V744,C159V1131,C159V1311,C159V1407:std_logic_vector(8 downto 0);
signal V187C160,V566C160,V623C160,V745C160,V1132C160,V1312C160,V1408C160,C160V187,C160V566,C160V623,C160V745,C160V1132,C160V1312,C160V1408:std_logic_vector(8 downto 0);
signal V188C161,V567C161,V624C161,V746C161,V1133C161,V1313C161,V1409C161,C161V188,C161V567,C161V624,C161V746,C161V1133,C161V1313,C161V1409:std_logic_vector(8 downto 0);
signal V189C162,V568C162,V625C162,V747C162,V1134C162,V1314C162,V1410C162,C162V189,C162V568,C162V625,C162V747,C162V1134,C162V1314,C162V1410:std_logic_vector(8 downto 0);
signal V190C163,V569C163,V626C163,V748C163,V1135C163,V1315C163,V1411C163,C163V190,C163V569,C163V626,C163V748,C163V1135,C163V1315,C163V1411:std_logic_vector(8 downto 0);
signal V191C164,V570C164,V627C164,V749C164,V1136C164,V1316C164,V1412C164,C164V191,C164V570,C164V627,C164V749,C164V1136,C164V1316,C164V1412:std_logic_vector(8 downto 0);
signal V192C165,V571C165,V628C165,V750C165,V1137C165,V1317C165,V1413C165,C165V192,C165V571,C165V628,C165V750,C165V1137,C165V1317,C165V1413:std_logic_vector(8 downto 0);
signal V97C166,V572C166,V629C166,V751C166,V1138C166,V1318C166,V1414C166,C166V97,C166V572,C166V629,C166V751,C166V1138,C166V1318,C166V1414:std_logic_vector(8 downto 0);
signal V98C167,V573C167,V630C167,V752C167,V1139C167,V1319C167,V1415C167,C167V98,C167V573,C167V630,C167V752,C167V1139,C167V1319,C167V1415:std_logic_vector(8 downto 0);
signal V99C168,V574C168,V631C168,V753C168,V1140C168,V1320C168,V1416C168,C168V99,C168V574,C168V631,C168V753,C168V1140,C168V1320,C168V1416:std_logic_vector(8 downto 0);
signal V100C169,V575C169,V632C169,V754C169,V1141C169,V1321C169,V1417C169,C169V100,C169V575,C169V632,C169V754,C169V1141,C169V1321,C169V1417:std_logic_vector(8 downto 0);
signal V101C170,V576C170,V633C170,V755C170,V1142C170,V1322C170,V1418C170,C170V101,C170V576,C170V633,C170V755,C170V1142,C170V1322,C170V1418:std_logic_vector(8 downto 0);
signal V102C171,V481C171,V634C171,V756C171,V1143C171,V1323C171,V1419C171,C171V102,C171V481,C171V634,C171V756,C171V1143,C171V1323,C171V1419:std_logic_vector(8 downto 0);
signal V103C172,V482C172,V635C172,V757C172,V1144C172,V1324C172,V1420C172,C172V103,C172V482,C172V635,C172V757,C172V1144,C172V1324,C172V1420:std_logic_vector(8 downto 0);
signal V104C173,V483C173,V636C173,V758C173,V1145C173,V1325C173,V1421C173,C173V104,C173V483,C173V636,C173V758,C173V1145,C173V1325,C173V1421:std_logic_vector(8 downto 0);
signal V105C174,V484C174,V637C174,V759C174,V1146C174,V1326C174,V1422C174,C174V105,C174V484,C174V637,C174V759,C174V1146,C174V1326,C174V1422:std_logic_vector(8 downto 0);
signal V106C175,V485C175,V638C175,V760C175,V1147C175,V1327C175,V1423C175,C175V106,C175V485,C175V638,C175V760,C175V1147,C175V1327,C175V1423:std_logic_vector(8 downto 0);
signal V107C176,V486C176,V639C176,V761C176,V1148C176,V1328C176,V1424C176,C176V107,C176V486,C176V639,C176V761,C176V1148,C176V1328,C176V1424:std_logic_vector(8 downto 0);
signal V108C177,V487C177,V640C177,V762C177,V1149C177,V1329C177,V1425C177,C177V108,C177V487,C177V640,C177V762,C177V1149,C177V1329,C177V1425:std_logic_vector(8 downto 0);
signal V109C178,V488C178,V641C178,V763C178,V1150C178,V1330C178,V1426C178,C178V109,C178V488,C178V641,C178V763,C178V1150,C178V1330,C178V1426:std_logic_vector(8 downto 0);
signal V110C179,V489C179,V642C179,V764C179,V1151C179,V1331C179,V1427C179,C179V110,C179V489,C179V642,C179V764,C179V1151,C179V1331,C179V1427:std_logic_vector(8 downto 0);
signal V111C180,V490C180,V643C180,V765C180,V1152C180,V1332C180,V1428C180,C180V111,C180V490,C180V643,C180V765,C180V1152,C180V1332,C180V1428:std_logic_vector(8 downto 0);
signal V112C181,V491C181,V644C181,V766C181,V1057C181,V1333C181,V1429C181,C181V112,C181V491,C181V644,C181V766,C181V1057,C181V1333,C181V1429:std_logic_vector(8 downto 0);
signal V113C182,V492C182,V645C182,V767C182,V1058C182,V1334C182,V1430C182,C182V113,C182V492,C182V645,C182V767,C182V1058,C182V1334,C182V1430:std_logic_vector(8 downto 0);
signal V114C183,V493C183,V646C183,V768C183,V1059C183,V1335C183,V1431C183,C183V114,C183V493,C183V646,C183V768,C183V1059,C183V1335,C183V1431:std_logic_vector(8 downto 0);
signal V115C184,V494C184,V647C184,V673C184,V1060C184,V1336C184,V1432C184,C184V115,C184V494,C184V647,C184V673,C184V1060,C184V1336,C184V1432:std_logic_vector(8 downto 0);
signal V116C185,V495C185,V648C185,V674C185,V1061C185,V1337C185,V1433C185,C185V116,C185V495,C185V648,C185V674,C185V1061,C185V1337,C185V1433:std_logic_vector(8 downto 0);
signal V117C186,V496C186,V649C186,V675C186,V1062C186,V1338C186,V1434C186,C186V117,C186V496,C186V649,C186V675,C186V1062,C186V1338,C186V1434:std_logic_vector(8 downto 0);
signal V118C187,V497C187,V650C187,V676C187,V1063C187,V1339C187,V1435C187,C187V118,C187V497,C187V650,C187V676,C187V1063,C187V1339,C187V1435:std_logic_vector(8 downto 0);
signal V119C188,V498C188,V651C188,V677C188,V1064C188,V1340C188,V1436C188,C188V119,C188V498,C188V651,C188V677,C188V1064,C188V1340,C188V1436:std_logic_vector(8 downto 0);
signal V120C189,V499C189,V652C189,V678C189,V1065C189,V1341C189,V1437C189,C189V120,C189V499,C189V652,C189V678,C189V1065,C189V1341,C189V1437:std_logic_vector(8 downto 0);
signal V121C190,V500C190,V653C190,V679C190,V1066C190,V1342C190,V1438C190,C190V121,C190V500,C190V653,C190V679,C190V1066,C190V1342,C190V1438:std_logic_vector(8 downto 0);
signal V122C191,V501C191,V654C191,V680C191,V1067C191,V1343C191,V1439C191,C191V122,C191V501,C191V654,C191V680,C191V1067,C191V1343,C191V1439:std_logic_vector(8 downto 0);
signal V123C192,V502C192,V655C192,V681C192,V1068C192,V1344C192,V1440C192,C192V123,C192V502,C192V655,C192V681,C192V1068,C192V1344,C192V1440:std_logic_vector(8 downto 0);
signal V313C193,V407C193,V562C193,V706C193,V1057C193,V1345C193,V1441C193,C193V313,C193V407,C193V562,C193V706,C193V1057,C193V1345,C193V1441:std_logic_vector(8 downto 0);
signal V314C194,V408C194,V563C194,V707C194,V1058C194,V1346C194,V1442C194,C194V314,C194V408,C194V563,C194V707,C194V1058,C194V1346,C194V1442:std_logic_vector(8 downto 0);
signal V315C195,V409C195,V564C195,V708C195,V1059C195,V1347C195,V1443C195,C195V315,C195V409,C195V564,C195V708,C195V1059,C195V1347,C195V1443:std_logic_vector(8 downto 0);
signal V316C196,V410C196,V565C196,V709C196,V1060C196,V1348C196,V1444C196,C196V316,C196V410,C196V565,C196V709,C196V1060,C196V1348,C196V1444:std_logic_vector(8 downto 0);
signal V317C197,V411C197,V566C197,V710C197,V1061C197,V1349C197,V1445C197,C197V317,C197V411,C197V566,C197V710,C197V1061,C197V1349,C197V1445:std_logic_vector(8 downto 0);
signal V318C198,V412C198,V567C198,V711C198,V1062C198,V1350C198,V1446C198,C198V318,C198V412,C198V567,C198V711,C198V1062,C198V1350,C198V1446:std_logic_vector(8 downto 0);
signal V319C199,V413C199,V568C199,V712C199,V1063C199,V1351C199,V1447C199,C199V319,C199V413,C199V568,C199V712,C199V1063,C199V1351,C199V1447:std_logic_vector(8 downto 0);
signal V320C200,V414C200,V569C200,V713C200,V1064C200,V1352C200,V1448C200,C200V320,C200V414,C200V569,C200V713,C200V1064,C200V1352,C200V1448:std_logic_vector(8 downto 0);
signal V321C201,V415C201,V570C201,V714C201,V1065C201,V1353C201,V1449C201,C201V321,C201V415,C201V570,C201V714,C201V1065,C201V1353,C201V1449:std_logic_vector(8 downto 0);
signal V322C202,V416C202,V571C202,V715C202,V1066C202,V1354C202,V1450C202,C202V322,C202V416,C202V571,C202V715,C202V1066,C202V1354,C202V1450:std_logic_vector(8 downto 0);
signal V323C203,V417C203,V572C203,V716C203,V1067C203,V1355C203,V1451C203,C203V323,C203V417,C203V572,C203V716,C203V1067,C203V1355,C203V1451:std_logic_vector(8 downto 0);
signal V324C204,V418C204,V573C204,V717C204,V1068C204,V1356C204,V1452C204,C204V324,C204V418,C204V573,C204V717,C204V1068,C204V1356,C204V1452:std_logic_vector(8 downto 0);
signal V325C205,V419C205,V574C205,V718C205,V1069C205,V1357C205,V1453C205,C205V325,C205V419,C205V574,C205V718,C205V1069,C205V1357,C205V1453:std_logic_vector(8 downto 0);
signal V326C206,V420C206,V575C206,V719C206,V1070C206,V1358C206,V1454C206,C206V326,C206V420,C206V575,C206V719,C206V1070,C206V1358,C206V1454:std_logic_vector(8 downto 0);
signal V327C207,V421C207,V576C207,V720C207,V1071C207,V1359C207,V1455C207,C207V327,C207V421,C207V576,C207V720,C207V1071,C207V1359,C207V1455:std_logic_vector(8 downto 0);
signal V328C208,V422C208,V481C208,V721C208,V1072C208,V1360C208,V1456C208,C208V328,C208V422,C208V481,C208V721,C208V1072,C208V1360,C208V1456:std_logic_vector(8 downto 0);
signal V329C209,V423C209,V482C209,V722C209,V1073C209,V1361C209,V1457C209,C209V329,C209V423,C209V482,C209V722,C209V1073,C209V1361,C209V1457:std_logic_vector(8 downto 0);
signal V330C210,V424C210,V483C210,V723C210,V1074C210,V1362C210,V1458C210,C210V330,C210V424,C210V483,C210V723,C210V1074,C210V1362,C210V1458:std_logic_vector(8 downto 0);
signal V331C211,V425C211,V484C211,V724C211,V1075C211,V1363C211,V1459C211,C211V331,C211V425,C211V484,C211V724,C211V1075,C211V1363,C211V1459:std_logic_vector(8 downto 0);
signal V332C212,V426C212,V485C212,V725C212,V1076C212,V1364C212,V1460C212,C212V332,C212V426,C212V485,C212V725,C212V1076,C212V1364,C212V1460:std_logic_vector(8 downto 0);
signal V333C213,V427C213,V486C213,V726C213,V1077C213,V1365C213,V1461C213,C213V333,C213V427,C213V486,C213V726,C213V1077,C213V1365,C213V1461:std_logic_vector(8 downto 0);
signal V334C214,V428C214,V487C214,V727C214,V1078C214,V1366C214,V1462C214,C214V334,C214V428,C214V487,C214V727,C214V1078,C214V1366,C214V1462:std_logic_vector(8 downto 0);
signal V335C215,V429C215,V488C215,V728C215,V1079C215,V1367C215,V1463C215,C215V335,C215V429,C215V488,C215V728,C215V1079,C215V1367,C215V1463:std_logic_vector(8 downto 0);
signal V336C216,V430C216,V489C216,V729C216,V1080C216,V1368C216,V1464C216,C216V336,C216V430,C216V489,C216V729,C216V1080,C216V1368,C216V1464:std_logic_vector(8 downto 0);
signal V337C217,V431C217,V490C217,V730C217,V1081C217,V1369C217,V1465C217,C217V337,C217V431,C217V490,C217V730,C217V1081,C217V1369,C217V1465:std_logic_vector(8 downto 0);
signal V338C218,V432C218,V491C218,V731C218,V1082C218,V1370C218,V1466C218,C218V338,C218V432,C218V491,C218V731,C218V1082,C218V1370,C218V1466:std_logic_vector(8 downto 0);
signal V339C219,V433C219,V492C219,V732C219,V1083C219,V1371C219,V1467C219,C219V339,C219V433,C219V492,C219V732,C219V1083,C219V1371,C219V1467:std_logic_vector(8 downto 0);
signal V340C220,V434C220,V493C220,V733C220,V1084C220,V1372C220,V1468C220,C220V340,C220V434,C220V493,C220V733,C220V1084,C220V1372,C220V1468:std_logic_vector(8 downto 0);
signal V341C221,V435C221,V494C221,V734C221,V1085C221,V1373C221,V1469C221,C221V341,C221V435,C221V494,C221V734,C221V1085,C221V1373,C221V1469:std_logic_vector(8 downto 0);
signal V342C222,V436C222,V495C222,V735C222,V1086C222,V1374C222,V1470C222,C222V342,C222V436,C222V495,C222V735,C222V1086,C222V1374,C222V1470:std_logic_vector(8 downto 0);
signal V343C223,V437C223,V496C223,V736C223,V1087C223,V1375C223,V1471C223,C223V343,C223V437,C223V496,C223V736,C223V1087,C223V1375,C223V1471:std_logic_vector(8 downto 0);
signal V344C224,V438C224,V497C224,V737C224,V1088C224,V1376C224,V1472C224,C224V344,C224V438,C224V497,C224V737,C224V1088,C224V1376,C224V1472:std_logic_vector(8 downto 0);
signal V345C225,V439C225,V498C225,V738C225,V1089C225,V1377C225,V1473C225,C225V345,C225V439,C225V498,C225V738,C225V1089,C225V1377,C225V1473:std_logic_vector(8 downto 0);
signal V346C226,V440C226,V499C226,V739C226,V1090C226,V1378C226,V1474C226,C226V346,C226V440,C226V499,C226V739,C226V1090,C226V1378,C226V1474:std_logic_vector(8 downto 0);
signal V347C227,V441C227,V500C227,V740C227,V1091C227,V1379C227,V1475C227,C227V347,C227V441,C227V500,C227V740,C227V1091,C227V1379,C227V1475:std_logic_vector(8 downto 0);
signal V348C228,V442C228,V501C228,V741C228,V1092C228,V1380C228,V1476C228,C228V348,C228V442,C228V501,C228V741,C228V1092,C228V1380,C228V1476:std_logic_vector(8 downto 0);
signal V349C229,V443C229,V502C229,V742C229,V1093C229,V1381C229,V1477C229,C229V349,C229V443,C229V502,C229V742,C229V1093,C229V1381,C229V1477:std_logic_vector(8 downto 0);
signal V350C230,V444C230,V503C230,V743C230,V1094C230,V1382C230,V1478C230,C230V350,C230V444,C230V503,C230V743,C230V1094,C230V1382,C230V1478:std_logic_vector(8 downto 0);
signal V351C231,V445C231,V504C231,V744C231,V1095C231,V1383C231,V1479C231,C231V351,C231V445,C231V504,C231V744,C231V1095,C231V1383,C231V1479:std_logic_vector(8 downto 0);
signal V352C232,V446C232,V505C232,V745C232,V1096C232,V1384C232,V1480C232,C232V352,C232V446,C232V505,C232V745,C232V1096,C232V1384,C232V1480:std_logic_vector(8 downto 0);
signal V353C233,V447C233,V506C233,V746C233,V1097C233,V1385C233,V1481C233,C233V353,C233V447,C233V506,C233V746,C233V1097,C233V1385,C233V1481:std_logic_vector(8 downto 0);
signal V354C234,V448C234,V507C234,V747C234,V1098C234,V1386C234,V1482C234,C234V354,C234V448,C234V507,C234V747,C234V1098,C234V1386,C234V1482:std_logic_vector(8 downto 0);
signal V355C235,V449C235,V508C235,V748C235,V1099C235,V1387C235,V1483C235,C235V355,C235V449,C235V508,C235V748,C235V1099,C235V1387,C235V1483:std_logic_vector(8 downto 0);
signal V356C236,V450C236,V509C236,V749C236,V1100C236,V1388C236,V1484C236,C236V356,C236V450,C236V509,C236V749,C236V1100,C236V1388,C236V1484:std_logic_vector(8 downto 0);
signal V357C237,V451C237,V510C237,V750C237,V1101C237,V1389C237,V1485C237,C237V357,C237V451,C237V510,C237V750,C237V1101,C237V1389,C237V1485:std_logic_vector(8 downto 0);
signal V358C238,V452C238,V511C238,V751C238,V1102C238,V1390C238,V1486C238,C238V358,C238V452,C238V511,C238V751,C238V1102,C238V1390,C238V1486:std_logic_vector(8 downto 0);
signal V359C239,V453C239,V512C239,V752C239,V1103C239,V1391C239,V1487C239,C239V359,C239V453,C239V512,C239V752,C239V1103,C239V1391,C239V1487:std_logic_vector(8 downto 0);
signal V360C240,V454C240,V513C240,V753C240,V1104C240,V1392C240,V1488C240,C240V360,C240V454,C240V513,C240V753,C240V1104,C240V1392,C240V1488:std_logic_vector(8 downto 0);
signal V361C241,V455C241,V514C241,V754C241,V1105C241,V1393C241,V1489C241,C241V361,C241V455,C241V514,C241V754,C241V1105,C241V1393,C241V1489:std_logic_vector(8 downto 0);
signal V362C242,V456C242,V515C242,V755C242,V1106C242,V1394C242,V1490C242,C242V362,C242V456,C242V515,C242V755,C242V1106,C242V1394,C242V1490:std_logic_vector(8 downto 0);
signal V363C243,V457C243,V516C243,V756C243,V1107C243,V1395C243,V1491C243,C243V363,C243V457,C243V516,C243V756,C243V1107,C243V1395,C243V1491:std_logic_vector(8 downto 0);
signal V364C244,V458C244,V517C244,V757C244,V1108C244,V1396C244,V1492C244,C244V364,C244V458,C244V517,C244V757,C244V1108,C244V1396,C244V1492:std_logic_vector(8 downto 0);
signal V365C245,V459C245,V518C245,V758C245,V1109C245,V1397C245,V1493C245,C245V365,C245V459,C245V518,C245V758,C245V1109,C245V1397,C245V1493:std_logic_vector(8 downto 0);
signal V366C246,V460C246,V519C246,V759C246,V1110C246,V1398C246,V1494C246,C246V366,C246V460,C246V519,C246V759,C246V1110,C246V1398,C246V1494:std_logic_vector(8 downto 0);
signal V367C247,V461C247,V520C247,V760C247,V1111C247,V1399C247,V1495C247,C247V367,C247V461,C247V520,C247V760,C247V1111,C247V1399,C247V1495:std_logic_vector(8 downto 0);
signal V368C248,V462C248,V521C248,V761C248,V1112C248,V1400C248,V1496C248,C248V368,C248V462,C248V521,C248V761,C248V1112,C248V1400,C248V1496:std_logic_vector(8 downto 0);
signal V369C249,V463C249,V522C249,V762C249,V1113C249,V1401C249,V1497C249,C249V369,C249V463,C249V522,C249V762,C249V1113,C249V1401,C249V1497:std_logic_vector(8 downto 0);
signal V370C250,V464C250,V523C250,V763C250,V1114C250,V1402C250,V1498C250,C250V370,C250V464,C250V523,C250V763,C250V1114,C250V1402,C250V1498:std_logic_vector(8 downto 0);
signal V371C251,V465C251,V524C251,V764C251,V1115C251,V1403C251,V1499C251,C251V371,C251V465,C251V524,C251V764,C251V1115,C251V1403,C251V1499:std_logic_vector(8 downto 0);
signal V372C252,V466C252,V525C252,V765C252,V1116C252,V1404C252,V1500C252,C252V372,C252V466,C252V525,C252V765,C252V1116,C252V1404,C252V1500:std_logic_vector(8 downto 0);
signal V373C253,V467C253,V526C253,V766C253,V1117C253,V1405C253,V1501C253,C253V373,C253V467,C253V526,C253V766,C253V1117,C253V1405,C253V1501:std_logic_vector(8 downto 0);
signal V374C254,V468C254,V527C254,V767C254,V1118C254,V1406C254,V1502C254,C254V374,C254V468,C254V527,C254V767,C254V1118,C254V1406,C254V1502:std_logic_vector(8 downto 0);
signal V375C255,V469C255,V528C255,V768C255,V1119C255,V1407C255,V1503C255,C255V375,C255V469,C255V528,C255V768,C255V1119,C255V1407,C255V1503:std_logic_vector(8 downto 0);
signal V376C256,V470C256,V529C256,V673C256,V1120C256,V1408C256,V1504C256,C256V376,C256V470,C256V529,C256V673,C256V1120,C256V1408,C256V1504:std_logic_vector(8 downto 0);
signal V377C257,V471C257,V530C257,V674C257,V1121C257,V1409C257,V1505C257,C257V377,C257V471,C257V530,C257V674,C257V1121,C257V1409,C257V1505:std_logic_vector(8 downto 0);
signal V378C258,V472C258,V531C258,V675C258,V1122C258,V1410C258,V1506C258,C258V378,C258V472,C258V531,C258V675,C258V1122,C258V1410,C258V1506:std_logic_vector(8 downto 0);
signal V379C259,V473C259,V532C259,V676C259,V1123C259,V1411C259,V1507C259,C259V379,C259V473,C259V532,C259V676,C259V1123,C259V1411,C259V1507:std_logic_vector(8 downto 0);
signal V380C260,V474C260,V533C260,V677C260,V1124C260,V1412C260,V1508C260,C260V380,C260V474,C260V533,C260V677,C260V1124,C260V1412,C260V1508:std_logic_vector(8 downto 0);
signal V381C261,V475C261,V534C261,V678C261,V1125C261,V1413C261,V1509C261,C261V381,C261V475,C261V534,C261V678,C261V1125,C261V1413,C261V1509:std_logic_vector(8 downto 0);
signal V382C262,V476C262,V535C262,V679C262,V1126C262,V1414C262,V1510C262,C262V382,C262V476,C262V535,C262V679,C262V1126,C262V1414,C262V1510:std_logic_vector(8 downto 0);
signal V383C263,V477C263,V536C263,V680C263,V1127C263,V1415C263,V1511C263,C263V383,C263V477,C263V536,C263V680,C263V1127,C263V1415,C263V1511:std_logic_vector(8 downto 0);
signal V384C264,V478C264,V537C264,V681C264,V1128C264,V1416C264,V1512C264,C264V384,C264V478,C264V537,C264V681,C264V1128,C264V1416,C264V1512:std_logic_vector(8 downto 0);
signal V289C265,V479C265,V538C265,V682C265,V1129C265,V1417C265,V1513C265,C265V289,C265V479,C265V538,C265V682,C265V1129,C265V1417,C265V1513:std_logic_vector(8 downto 0);
signal V290C266,V480C266,V539C266,V683C266,V1130C266,V1418C266,V1514C266,C266V290,C266V480,C266V539,C266V683,C266V1130,C266V1418,C266V1514:std_logic_vector(8 downto 0);
signal V291C267,V385C267,V540C267,V684C267,V1131C267,V1419C267,V1515C267,C267V291,C267V385,C267V540,C267V684,C267V1131,C267V1419,C267V1515:std_logic_vector(8 downto 0);
signal V292C268,V386C268,V541C268,V685C268,V1132C268,V1420C268,V1516C268,C268V292,C268V386,C268V541,C268V685,C268V1132,C268V1420,C268V1516:std_logic_vector(8 downto 0);
signal V293C269,V387C269,V542C269,V686C269,V1133C269,V1421C269,V1517C269,C269V293,C269V387,C269V542,C269V686,C269V1133,C269V1421,C269V1517:std_logic_vector(8 downto 0);
signal V294C270,V388C270,V543C270,V687C270,V1134C270,V1422C270,V1518C270,C270V294,C270V388,C270V543,C270V687,C270V1134,C270V1422,C270V1518:std_logic_vector(8 downto 0);
signal V295C271,V389C271,V544C271,V688C271,V1135C271,V1423C271,V1519C271,C271V295,C271V389,C271V544,C271V688,C271V1135,C271V1423,C271V1519:std_logic_vector(8 downto 0);
signal V296C272,V390C272,V545C272,V689C272,V1136C272,V1424C272,V1520C272,C272V296,C272V390,C272V545,C272V689,C272V1136,C272V1424,C272V1520:std_logic_vector(8 downto 0);
signal V297C273,V391C273,V546C273,V690C273,V1137C273,V1425C273,V1521C273,C273V297,C273V391,C273V546,C273V690,C273V1137,C273V1425,C273V1521:std_logic_vector(8 downto 0);
signal V298C274,V392C274,V547C274,V691C274,V1138C274,V1426C274,V1522C274,C274V298,C274V392,C274V547,C274V691,C274V1138,C274V1426,C274V1522:std_logic_vector(8 downto 0);
signal V299C275,V393C275,V548C275,V692C275,V1139C275,V1427C275,V1523C275,C275V299,C275V393,C275V548,C275V692,C275V1139,C275V1427,C275V1523:std_logic_vector(8 downto 0);
signal V300C276,V394C276,V549C276,V693C276,V1140C276,V1428C276,V1524C276,C276V300,C276V394,C276V549,C276V693,C276V1140,C276V1428,C276V1524:std_logic_vector(8 downto 0);
signal V301C277,V395C277,V550C277,V694C277,V1141C277,V1429C277,V1525C277,C277V301,C277V395,C277V550,C277V694,C277V1141,C277V1429,C277V1525:std_logic_vector(8 downto 0);
signal V302C278,V396C278,V551C278,V695C278,V1142C278,V1430C278,V1526C278,C278V302,C278V396,C278V551,C278V695,C278V1142,C278V1430,C278V1526:std_logic_vector(8 downto 0);
signal V303C279,V397C279,V552C279,V696C279,V1143C279,V1431C279,V1527C279,C279V303,C279V397,C279V552,C279V696,C279V1143,C279V1431,C279V1527:std_logic_vector(8 downto 0);
signal V304C280,V398C280,V553C280,V697C280,V1144C280,V1432C280,V1528C280,C280V304,C280V398,C280V553,C280V697,C280V1144,C280V1432,C280V1528:std_logic_vector(8 downto 0);
signal V305C281,V399C281,V554C281,V698C281,V1145C281,V1433C281,V1529C281,C281V305,C281V399,C281V554,C281V698,C281V1145,C281V1433,C281V1529:std_logic_vector(8 downto 0);
signal V306C282,V400C282,V555C282,V699C282,V1146C282,V1434C282,V1530C282,C282V306,C282V400,C282V555,C282V699,C282V1146,C282V1434,C282V1530:std_logic_vector(8 downto 0);
signal V307C283,V401C283,V556C283,V700C283,V1147C283,V1435C283,V1531C283,C283V307,C283V401,C283V556,C283V700,C283V1147,C283V1435,C283V1531:std_logic_vector(8 downto 0);
signal V308C284,V402C284,V557C284,V701C284,V1148C284,V1436C284,V1532C284,C284V308,C284V402,C284V557,C284V701,C284V1148,C284V1436,C284V1532:std_logic_vector(8 downto 0);
signal V309C285,V403C285,V558C285,V702C285,V1149C285,V1437C285,V1533C285,C285V309,C285V403,C285V558,C285V702,C285V1149,C285V1437,C285V1533:std_logic_vector(8 downto 0);
signal V310C286,V404C286,V559C286,V703C286,V1150C286,V1438C286,V1534C286,C286V310,C286V404,C286V559,C286V703,C286V1150,C286V1438,C286V1534:std_logic_vector(8 downto 0);
signal V311C287,V405C287,V560C287,V704C287,V1151C287,V1439C287,V1535C287,C287V311,C287V405,C287V560,C287V704,C287V1151,C287V1439,C287V1535:std_logic_vector(8 downto 0);
signal V312C288,V406C288,V561C288,V705C288,V1152C288,V1440C288,V1536C288,C288V312,C288V406,C288V561,C288V705,C288V1152,C288V1440,C288V1536:std_logic_vector(8 downto 0);
signal V62C289,V240C289,V834C289,V890C289,V1441C289,V1537C289,C289V62,C289V240,C289V834,C289V890,C289V1441,C289V1537:std_logic_vector(8 downto 0);
signal V63C290,V241C290,V835C290,V891C290,V1442C290,V1538C290,C290V63,C290V241,C290V835,C290V891,C290V1442,C290V1538:std_logic_vector(8 downto 0);
signal V64C291,V242C291,V836C291,V892C291,V1443C291,V1539C291,C291V64,C291V242,C291V836,C291V892,C291V1443,C291V1539:std_logic_vector(8 downto 0);
signal V65C292,V243C292,V837C292,V893C292,V1444C292,V1540C292,C292V65,C292V243,C292V837,C292V893,C292V1444,C292V1540:std_logic_vector(8 downto 0);
signal V66C293,V244C293,V838C293,V894C293,V1445C293,V1541C293,C293V66,C293V244,C293V838,C293V894,C293V1445,C293V1541:std_logic_vector(8 downto 0);
signal V67C294,V245C294,V839C294,V895C294,V1446C294,V1542C294,C294V67,C294V245,C294V839,C294V895,C294V1446,C294V1542:std_logic_vector(8 downto 0);
signal V68C295,V246C295,V840C295,V896C295,V1447C295,V1543C295,C295V68,C295V246,C295V840,C295V896,C295V1447,C295V1543:std_logic_vector(8 downto 0);
signal V69C296,V247C296,V841C296,V897C296,V1448C296,V1544C296,C296V69,C296V247,C296V841,C296V897,C296V1448,C296V1544:std_logic_vector(8 downto 0);
signal V70C297,V248C297,V842C297,V898C297,V1449C297,V1545C297,C297V70,C297V248,C297V842,C297V898,C297V1449,C297V1545:std_logic_vector(8 downto 0);
signal V71C298,V249C298,V843C298,V899C298,V1450C298,V1546C298,C298V71,C298V249,C298V843,C298V899,C298V1450,C298V1546:std_logic_vector(8 downto 0);
signal V72C299,V250C299,V844C299,V900C299,V1451C299,V1547C299,C299V72,C299V250,C299V844,C299V900,C299V1451,C299V1547:std_logic_vector(8 downto 0);
signal V73C300,V251C300,V845C300,V901C300,V1452C300,V1548C300,C300V73,C300V251,C300V845,C300V901,C300V1452,C300V1548:std_logic_vector(8 downto 0);
signal V74C301,V252C301,V846C301,V902C301,V1453C301,V1549C301,C301V74,C301V252,C301V846,C301V902,C301V1453,C301V1549:std_logic_vector(8 downto 0);
signal V75C302,V253C302,V847C302,V903C302,V1454C302,V1550C302,C302V75,C302V253,C302V847,C302V903,C302V1454,C302V1550:std_logic_vector(8 downto 0);
signal V76C303,V254C303,V848C303,V904C303,V1455C303,V1551C303,C303V76,C303V254,C303V848,C303V904,C303V1455,C303V1551:std_logic_vector(8 downto 0);
signal V77C304,V255C304,V849C304,V905C304,V1456C304,V1552C304,C304V77,C304V255,C304V849,C304V905,C304V1456,C304V1552:std_logic_vector(8 downto 0);
signal V78C305,V256C305,V850C305,V906C305,V1457C305,V1553C305,C305V78,C305V256,C305V850,C305V906,C305V1457,C305V1553:std_logic_vector(8 downto 0);
signal V79C306,V257C306,V851C306,V907C306,V1458C306,V1554C306,C306V79,C306V257,C306V851,C306V907,C306V1458,C306V1554:std_logic_vector(8 downto 0);
signal V80C307,V258C307,V852C307,V908C307,V1459C307,V1555C307,C307V80,C307V258,C307V852,C307V908,C307V1459,C307V1555:std_logic_vector(8 downto 0);
signal V81C308,V259C308,V853C308,V909C308,V1460C308,V1556C308,C308V81,C308V259,C308V853,C308V909,C308V1460,C308V1556:std_logic_vector(8 downto 0);
signal V82C309,V260C309,V854C309,V910C309,V1461C309,V1557C309,C309V82,C309V260,C309V854,C309V910,C309V1461,C309V1557:std_logic_vector(8 downto 0);
signal V83C310,V261C310,V855C310,V911C310,V1462C310,V1558C310,C310V83,C310V261,C310V855,C310V911,C310V1462,C310V1558:std_logic_vector(8 downto 0);
signal V84C311,V262C311,V856C311,V912C311,V1463C311,V1559C311,C311V84,C311V262,C311V856,C311V912,C311V1463,C311V1559:std_logic_vector(8 downto 0);
signal V85C312,V263C312,V857C312,V913C312,V1464C312,V1560C312,C312V85,C312V263,C312V857,C312V913,C312V1464,C312V1560:std_logic_vector(8 downto 0);
signal V86C313,V264C313,V858C313,V914C313,V1465C313,V1561C313,C313V86,C313V264,C313V858,C313V914,C313V1465,C313V1561:std_logic_vector(8 downto 0);
signal V87C314,V265C314,V859C314,V915C314,V1466C314,V1562C314,C314V87,C314V265,C314V859,C314V915,C314V1466,C314V1562:std_logic_vector(8 downto 0);
signal V88C315,V266C315,V860C315,V916C315,V1467C315,V1563C315,C315V88,C315V266,C315V860,C315V916,C315V1467,C315V1563:std_logic_vector(8 downto 0);
signal V89C316,V267C316,V861C316,V917C316,V1468C316,V1564C316,C316V89,C316V267,C316V861,C316V917,C316V1468,C316V1564:std_logic_vector(8 downto 0);
signal V90C317,V268C317,V862C317,V918C317,V1469C317,V1565C317,C317V90,C317V268,C317V862,C317V918,C317V1469,C317V1565:std_logic_vector(8 downto 0);
signal V91C318,V269C318,V863C318,V919C318,V1470C318,V1566C318,C318V91,C318V269,C318V863,C318V919,C318V1470,C318V1566:std_logic_vector(8 downto 0);
signal V92C319,V270C319,V864C319,V920C319,V1471C319,V1567C319,C319V92,C319V270,C319V864,C319V920,C319V1471,C319V1567:std_logic_vector(8 downto 0);
signal V93C320,V271C320,V769C320,V921C320,V1472C320,V1568C320,C320V93,C320V271,C320V769,C320V921,C320V1472,C320V1568:std_logic_vector(8 downto 0);
signal V94C321,V272C321,V770C321,V922C321,V1473C321,V1569C321,C321V94,C321V272,C321V770,C321V922,C321V1473,C321V1569:std_logic_vector(8 downto 0);
signal V95C322,V273C322,V771C322,V923C322,V1474C322,V1570C322,C322V95,C322V273,C322V771,C322V923,C322V1474,C322V1570:std_logic_vector(8 downto 0);
signal V96C323,V274C323,V772C323,V924C323,V1475C323,V1571C323,C323V96,C323V274,C323V772,C323V924,C323V1475,C323V1571:std_logic_vector(8 downto 0);
signal V1C324,V275C324,V773C324,V925C324,V1476C324,V1572C324,C324V1,C324V275,C324V773,C324V925,C324V1476,C324V1572:std_logic_vector(8 downto 0);
signal V2C325,V276C325,V774C325,V926C325,V1477C325,V1573C325,C325V2,C325V276,C325V774,C325V926,C325V1477,C325V1573:std_logic_vector(8 downto 0);
signal V3C326,V277C326,V775C326,V927C326,V1478C326,V1574C326,C326V3,C326V277,C326V775,C326V927,C326V1478,C326V1574:std_logic_vector(8 downto 0);
signal V4C327,V278C327,V776C327,V928C327,V1479C327,V1575C327,C327V4,C327V278,C327V776,C327V928,C327V1479,C327V1575:std_logic_vector(8 downto 0);
signal V5C328,V279C328,V777C328,V929C328,V1480C328,V1576C328,C328V5,C328V279,C328V777,C328V929,C328V1480,C328V1576:std_logic_vector(8 downto 0);
signal V6C329,V280C329,V778C329,V930C329,V1481C329,V1577C329,C329V6,C329V280,C329V778,C329V930,C329V1481,C329V1577:std_logic_vector(8 downto 0);
signal V7C330,V281C330,V779C330,V931C330,V1482C330,V1578C330,C330V7,C330V281,C330V779,C330V931,C330V1482,C330V1578:std_logic_vector(8 downto 0);
signal V8C331,V282C331,V780C331,V932C331,V1483C331,V1579C331,C331V8,C331V282,C331V780,C331V932,C331V1483,C331V1579:std_logic_vector(8 downto 0);
signal V9C332,V283C332,V781C332,V933C332,V1484C332,V1580C332,C332V9,C332V283,C332V781,C332V933,C332V1484,C332V1580:std_logic_vector(8 downto 0);
signal V10C333,V284C333,V782C333,V934C333,V1485C333,V1581C333,C333V10,C333V284,C333V782,C333V934,C333V1485,C333V1581:std_logic_vector(8 downto 0);
signal V11C334,V285C334,V783C334,V935C334,V1486C334,V1582C334,C334V11,C334V285,C334V783,C334V935,C334V1486,C334V1582:std_logic_vector(8 downto 0);
signal V12C335,V286C335,V784C335,V936C335,V1487C335,V1583C335,C335V12,C335V286,C335V784,C335V936,C335V1487,C335V1583:std_logic_vector(8 downto 0);
signal V13C336,V287C336,V785C336,V937C336,V1488C336,V1584C336,C336V13,C336V287,C336V785,C336V937,C336V1488,C336V1584:std_logic_vector(8 downto 0);
signal V14C337,V288C337,V786C337,V938C337,V1489C337,V1585C337,C337V14,C337V288,C337V786,C337V938,C337V1489,C337V1585:std_logic_vector(8 downto 0);
signal V15C338,V193C338,V787C338,V939C338,V1490C338,V1586C338,C338V15,C338V193,C338V787,C338V939,C338V1490,C338V1586:std_logic_vector(8 downto 0);
signal V16C339,V194C339,V788C339,V940C339,V1491C339,V1587C339,C339V16,C339V194,C339V788,C339V940,C339V1491,C339V1587:std_logic_vector(8 downto 0);
signal V17C340,V195C340,V789C340,V941C340,V1492C340,V1588C340,C340V17,C340V195,C340V789,C340V941,C340V1492,C340V1588:std_logic_vector(8 downto 0);
signal V18C341,V196C341,V790C341,V942C341,V1493C341,V1589C341,C341V18,C341V196,C341V790,C341V942,C341V1493,C341V1589:std_logic_vector(8 downto 0);
signal V19C342,V197C342,V791C342,V943C342,V1494C342,V1590C342,C342V19,C342V197,C342V791,C342V943,C342V1494,C342V1590:std_logic_vector(8 downto 0);
signal V20C343,V198C343,V792C343,V944C343,V1495C343,V1591C343,C343V20,C343V198,C343V792,C343V944,C343V1495,C343V1591:std_logic_vector(8 downto 0);
signal V21C344,V199C344,V793C344,V945C344,V1496C344,V1592C344,C344V21,C344V199,C344V793,C344V945,C344V1496,C344V1592:std_logic_vector(8 downto 0);
signal V22C345,V200C345,V794C345,V946C345,V1497C345,V1593C345,C345V22,C345V200,C345V794,C345V946,C345V1497,C345V1593:std_logic_vector(8 downto 0);
signal V23C346,V201C346,V795C346,V947C346,V1498C346,V1594C346,C346V23,C346V201,C346V795,C346V947,C346V1498,C346V1594:std_logic_vector(8 downto 0);
signal V24C347,V202C347,V796C347,V948C347,V1499C347,V1595C347,C347V24,C347V202,C347V796,C347V948,C347V1499,C347V1595:std_logic_vector(8 downto 0);
signal V25C348,V203C348,V797C348,V949C348,V1500C348,V1596C348,C348V25,C348V203,C348V797,C348V949,C348V1500,C348V1596:std_logic_vector(8 downto 0);
signal V26C349,V204C349,V798C349,V950C349,V1501C349,V1597C349,C349V26,C349V204,C349V798,C349V950,C349V1501,C349V1597:std_logic_vector(8 downto 0);
signal V27C350,V205C350,V799C350,V951C350,V1502C350,V1598C350,C350V27,C350V205,C350V799,C350V951,C350V1502,C350V1598:std_logic_vector(8 downto 0);
signal V28C351,V206C351,V800C351,V952C351,V1503C351,V1599C351,C351V28,C351V206,C351V800,C351V952,C351V1503,C351V1599:std_logic_vector(8 downto 0);
signal V29C352,V207C352,V801C352,V953C352,V1504C352,V1600C352,C352V29,C352V207,C352V801,C352V953,C352V1504,C352V1600:std_logic_vector(8 downto 0);
signal V30C353,V208C353,V802C353,V954C353,V1505C353,V1601C353,C353V30,C353V208,C353V802,C353V954,C353V1505,C353V1601:std_logic_vector(8 downto 0);
signal V31C354,V209C354,V803C354,V955C354,V1506C354,V1602C354,C354V31,C354V209,C354V803,C354V955,C354V1506,C354V1602:std_logic_vector(8 downto 0);
signal V32C355,V210C355,V804C355,V956C355,V1507C355,V1603C355,C355V32,C355V210,C355V804,C355V956,C355V1507,C355V1603:std_logic_vector(8 downto 0);
signal V33C356,V211C356,V805C356,V957C356,V1508C356,V1604C356,C356V33,C356V211,C356V805,C356V957,C356V1508,C356V1604:std_logic_vector(8 downto 0);
signal V34C357,V212C357,V806C357,V958C357,V1509C357,V1605C357,C357V34,C357V212,C357V806,C357V958,C357V1509,C357V1605:std_logic_vector(8 downto 0);
signal V35C358,V213C358,V807C358,V959C358,V1510C358,V1606C358,C358V35,C358V213,C358V807,C358V959,C358V1510,C358V1606:std_logic_vector(8 downto 0);
signal V36C359,V214C359,V808C359,V960C359,V1511C359,V1607C359,C359V36,C359V214,C359V808,C359V960,C359V1511,C359V1607:std_logic_vector(8 downto 0);
signal V37C360,V215C360,V809C360,V865C360,V1512C360,V1608C360,C360V37,C360V215,C360V809,C360V865,C360V1512,C360V1608:std_logic_vector(8 downto 0);
signal V38C361,V216C361,V810C361,V866C361,V1513C361,V1609C361,C361V38,C361V216,C361V810,C361V866,C361V1513,C361V1609:std_logic_vector(8 downto 0);
signal V39C362,V217C362,V811C362,V867C362,V1514C362,V1610C362,C362V39,C362V217,C362V811,C362V867,C362V1514,C362V1610:std_logic_vector(8 downto 0);
signal V40C363,V218C363,V812C363,V868C363,V1515C363,V1611C363,C363V40,C363V218,C363V812,C363V868,C363V1515,C363V1611:std_logic_vector(8 downto 0);
signal V41C364,V219C364,V813C364,V869C364,V1516C364,V1612C364,C364V41,C364V219,C364V813,C364V869,C364V1516,C364V1612:std_logic_vector(8 downto 0);
signal V42C365,V220C365,V814C365,V870C365,V1517C365,V1613C365,C365V42,C365V220,C365V814,C365V870,C365V1517,C365V1613:std_logic_vector(8 downto 0);
signal V43C366,V221C366,V815C366,V871C366,V1518C366,V1614C366,C366V43,C366V221,C366V815,C366V871,C366V1518,C366V1614:std_logic_vector(8 downto 0);
signal V44C367,V222C367,V816C367,V872C367,V1519C367,V1615C367,C367V44,C367V222,C367V816,C367V872,C367V1519,C367V1615:std_logic_vector(8 downto 0);
signal V45C368,V223C368,V817C368,V873C368,V1520C368,V1616C368,C368V45,C368V223,C368V817,C368V873,C368V1520,C368V1616:std_logic_vector(8 downto 0);
signal V46C369,V224C369,V818C369,V874C369,V1521C369,V1617C369,C369V46,C369V224,C369V818,C369V874,C369V1521,C369V1617:std_logic_vector(8 downto 0);
signal V47C370,V225C370,V819C370,V875C370,V1522C370,V1618C370,C370V47,C370V225,C370V819,C370V875,C370V1522,C370V1618:std_logic_vector(8 downto 0);
signal V48C371,V226C371,V820C371,V876C371,V1523C371,V1619C371,C371V48,C371V226,C371V820,C371V876,C371V1523,C371V1619:std_logic_vector(8 downto 0);
signal V49C372,V227C372,V821C372,V877C372,V1524C372,V1620C372,C372V49,C372V227,C372V821,C372V877,C372V1524,C372V1620:std_logic_vector(8 downto 0);
signal V50C373,V228C373,V822C373,V878C373,V1525C373,V1621C373,C373V50,C373V228,C373V822,C373V878,C373V1525,C373V1621:std_logic_vector(8 downto 0);
signal V51C374,V229C374,V823C374,V879C374,V1526C374,V1622C374,C374V51,C374V229,C374V823,C374V879,C374V1526,C374V1622:std_logic_vector(8 downto 0);
signal V52C375,V230C375,V824C375,V880C375,V1527C375,V1623C375,C375V52,C375V230,C375V824,C375V880,C375V1527,C375V1623:std_logic_vector(8 downto 0);
signal V53C376,V231C376,V825C376,V881C376,V1528C376,V1624C376,C376V53,C376V231,C376V825,C376V881,C376V1528,C376V1624:std_logic_vector(8 downto 0);
signal V54C377,V232C377,V826C377,V882C377,V1529C377,V1625C377,C377V54,C377V232,C377V826,C377V882,C377V1529,C377V1625:std_logic_vector(8 downto 0);
signal V55C378,V233C378,V827C378,V883C378,V1530C378,V1626C378,C378V55,C378V233,C378V827,C378V883,C378V1530,C378V1626:std_logic_vector(8 downto 0);
signal V56C379,V234C379,V828C379,V884C379,V1531C379,V1627C379,C379V56,C379V234,C379V828,C379V884,C379V1531,C379V1627:std_logic_vector(8 downto 0);
signal V57C380,V235C380,V829C380,V885C380,V1532C380,V1628C380,C380V57,C380V235,C380V829,C380V885,C380V1532,C380V1628:std_logic_vector(8 downto 0);
signal V58C381,V236C381,V830C381,V886C381,V1533C381,V1629C381,C381V58,C381V236,C381V830,C381V886,C381V1533,C381V1629:std_logic_vector(8 downto 0);
signal V59C382,V237C382,V831C382,V887C382,V1534C382,V1630C382,C382V59,C382V237,C382V831,C382V887,C382V1534,C382V1630:std_logic_vector(8 downto 0);
signal V60C383,V238C383,V832C383,V888C383,V1535C383,V1631C383,C383V60,C383V238,C383V832,C383V888,C383V1535,C383V1631:std_logic_vector(8 downto 0);
signal V61C384,V239C384,V833C384,V889C384,V1536C384,V1632C384,C384V61,C384V239,C384V833,C384V889,C384V1536,C384V1632:std_logic_vector(8 downto 0);
signal V232C385,V661C385,V906C385,V1033C385,V1537C385,V1633C385,C385V232,C385V661,C385V906,C385V1033,C385V1537,C385V1633:std_logic_vector(8 downto 0);
signal V233C386,V662C386,V907C386,V1034C386,V1538C386,V1634C386,C386V233,C386V662,C386V907,C386V1034,C386V1538,C386V1634:std_logic_vector(8 downto 0);
signal V234C387,V663C387,V908C387,V1035C387,V1539C387,V1635C387,C387V234,C387V663,C387V908,C387V1035,C387V1539,C387V1635:std_logic_vector(8 downto 0);
signal V235C388,V664C388,V909C388,V1036C388,V1540C388,V1636C388,C388V235,C388V664,C388V909,C388V1036,C388V1540,C388V1636:std_logic_vector(8 downto 0);
signal V236C389,V665C389,V910C389,V1037C389,V1541C389,V1637C389,C389V236,C389V665,C389V910,C389V1037,C389V1541,C389V1637:std_logic_vector(8 downto 0);
signal V237C390,V666C390,V911C390,V1038C390,V1542C390,V1638C390,C390V237,C390V666,C390V911,C390V1038,C390V1542,C390V1638:std_logic_vector(8 downto 0);
signal V238C391,V667C391,V912C391,V1039C391,V1543C391,V1639C391,C391V238,C391V667,C391V912,C391V1039,C391V1543,C391V1639:std_logic_vector(8 downto 0);
signal V239C392,V668C392,V913C392,V1040C392,V1544C392,V1640C392,C392V239,C392V668,C392V913,C392V1040,C392V1544,C392V1640:std_logic_vector(8 downto 0);
signal V240C393,V669C393,V914C393,V1041C393,V1545C393,V1641C393,C393V240,C393V669,C393V914,C393V1041,C393V1545,C393V1641:std_logic_vector(8 downto 0);
signal V241C394,V670C394,V915C394,V1042C394,V1546C394,V1642C394,C394V241,C394V670,C394V915,C394V1042,C394V1546,C394V1642:std_logic_vector(8 downto 0);
signal V242C395,V671C395,V916C395,V1043C395,V1547C395,V1643C395,C395V242,C395V671,C395V916,C395V1043,C395V1547,C395V1643:std_logic_vector(8 downto 0);
signal V243C396,V672C396,V917C396,V1044C396,V1548C396,V1644C396,C396V243,C396V672,C396V917,C396V1044,C396V1548,C396V1644:std_logic_vector(8 downto 0);
signal V244C397,V577C397,V918C397,V1045C397,V1549C397,V1645C397,C397V244,C397V577,C397V918,C397V1045,C397V1549,C397V1645:std_logic_vector(8 downto 0);
signal V245C398,V578C398,V919C398,V1046C398,V1550C398,V1646C398,C398V245,C398V578,C398V919,C398V1046,C398V1550,C398V1646:std_logic_vector(8 downto 0);
signal V246C399,V579C399,V920C399,V1047C399,V1551C399,V1647C399,C399V246,C399V579,C399V920,C399V1047,C399V1551,C399V1647:std_logic_vector(8 downto 0);
signal V247C400,V580C400,V921C400,V1048C400,V1552C400,V1648C400,C400V247,C400V580,C400V921,C400V1048,C400V1552,C400V1648:std_logic_vector(8 downto 0);
signal V248C401,V581C401,V922C401,V1049C401,V1553C401,V1649C401,C401V248,C401V581,C401V922,C401V1049,C401V1553,C401V1649:std_logic_vector(8 downto 0);
signal V249C402,V582C402,V923C402,V1050C402,V1554C402,V1650C402,C402V249,C402V582,C402V923,C402V1050,C402V1554,C402V1650:std_logic_vector(8 downto 0);
signal V250C403,V583C403,V924C403,V1051C403,V1555C403,V1651C403,C403V250,C403V583,C403V924,C403V1051,C403V1555,C403V1651:std_logic_vector(8 downto 0);
signal V251C404,V584C404,V925C404,V1052C404,V1556C404,V1652C404,C404V251,C404V584,C404V925,C404V1052,C404V1556,C404V1652:std_logic_vector(8 downto 0);
signal V252C405,V585C405,V926C405,V1053C405,V1557C405,V1653C405,C405V252,C405V585,C405V926,C405V1053,C405V1557,C405V1653:std_logic_vector(8 downto 0);
signal V253C406,V586C406,V927C406,V1054C406,V1558C406,V1654C406,C406V253,C406V586,C406V927,C406V1054,C406V1558,C406V1654:std_logic_vector(8 downto 0);
signal V254C407,V587C407,V928C407,V1055C407,V1559C407,V1655C407,C407V254,C407V587,C407V928,C407V1055,C407V1559,C407V1655:std_logic_vector(8 downto 0);
signal V255C408,V588C408,V929C408,V1056C408,V1560C408,V1656C408,C408V255,C408V588,C408V929,C408V1056,C408V1560,C408V1656:std_logic_vector(8 downto 0);
signal V256C409,V589C409,V930C409,V961C409,V1561C409,V1657C409,C409V256,C409V589,C409V930,C409V961,C409V1561,C409V1657:std_logic_vector(8 downto 0);
signal V257C410,V590C410,V931C410,V962C410,V1562C410,V1658C410,C410V257,C410V590,C410V931,C410V962,C410V1562,C410V1658:std_logic_vector(8 downto 0);
signal V258C411,V591C411,V932C411,V963C411,V1563C411,V1659C411,C411V258,C411V591,C411V932,C411V963,C411V1563,C411V1659:std_logic_vector(8 downto 0);
signal V259C412,V592C412,V933C412,V964C412,V1564C412,V1660C412,C412V259,C412V592,C412V933,C412V964,C412V1564,C412V1660:std_logic_vector(8 downto 0);
signal V260C413,V593C413,V934C413,V965C413,V1565C413,V1661C413,C413V260,C413V593,C413V934,C413V965,C413V1565,C413V1661:std_logic_vector(8 downto 0);
signal V261C414,V594C414,V935C414,V966C414,V1566C414,V1662C414,C414V261,C414V594,C414V935,C414V966,C414V1566,C414V1662:std_logic_vector(8 downto 0);
signal V262C415,V595C415,V936C415,V967C415,V1567C415,V1663C415,C415V262,C415V595,C415V936,C415V967,C415V1567,C415V1663:std_logic_vector(8 downto 0);
signal V263C416,V596C416,V937C416,V968C416,V1568C416,V1664C416,C416V263,C416V596,C416V937,C416V968,C416V1568,C416V1664:std_logic_vector(8 downto 0);
signal V264C417,V597C417,V938C417,V969C417,V1569C417,V1665C417,C417V264,C417V597,C417V938,C417V969,C417V1569,C417V1665:std_logic_vector(8 downto 0);
signal V265C418,V598C418,V939C418,V970C418,V1570C418,V1666C418,C418V265,C418V598,C418V939,C418V970,C418V1570,C418V1666:std_logic_vector(8 downto 0);
signal V266C419,V599C419,V940C419,V971C419,V1571C419,V1667C419,C419V266,C419V599,C419V940,C419V971,C419V1571,C419V1667:std_logic_vector(8 downto 0);
signal V267C420,V600C420,V941C420,V972C420,V1572C420,V1668C420,C420V267,C420V600,C420V941,C420V972,C420V1572,C420V1668:std_logic_vector(8 downto 0);
signal V268C421,V601C421,V942C421,V973C421,V1573C421,V1669C421,C421V268,C421V601,C421V942,C421V973,C421V1573,C421V1669:std_logic_vector(8 downto 0);
signal V269C422,V602C422,V943C422,V974C422,V1574C422,V1670C422,C422V269,C422V602,C422V943,C422V974,C422V1574,C422V1670:std_logic_vector(8 downto 0);
signal V270C423,V603C423,V944C423,V975C423,V1575C423,V1671C423,C423V270,C423V603,C423V944,C423V975,C423V1575,C423V1671:std_logic_vector(8 downto 0);
signal V271C424,V604C424,V945C424,V976C424,V1576C424,V1672C424,C424V271,C424V604,C424V945,C424V976,C424V1576,C424V1672:std_logic_vector(8 downto 0);
signal V272C425,V605C425,V946C425,V977C425,V1577C425,V1673C425,C425V272,C425V605,C425V946,C425V977,C425V1577,C425V1673:std_logic_vector(8 downto 0);
signal V273C426,V606C426,V947C426,V978C426,V1578C426,V1674C426,C426V273,C426V606,C426V947,C426V978,C426V1578,C426V1674:std_logic_vector(8 downto 0);
signal V274C427,V607C427,V948C427,V979C427,V1579C427,V1675C427,C427V274,C427V607,C427V948,C427V979,C427V1579,C427V1675:std_logic_vector(8 downto 0);
signal V275C428,V608C428,V949C428,V980C428,V1580C428,V1676C428,C428V275,C428V608,C428V949,C428V980,C428V1580,C428V1676:std_logic_vector(8 downto 0);
signal V276C429,V609C429,V950C429,V981C429,V1581C429,V1677C429,C429V276,C429V609,C429V950,C429V981,C429V1581,C429V1677:std_logic_vector(8 downto 0);
signal V277C430,V610C430,V951C430,V982C430,V1582C430,V1678C430,C430V277,C430V610,C430V951,C430V982,C430V1582,C430V1678:std_logic_vector(8 downto 0);
signal V278C431,V611C431,V952C431,V983C431,V1583C431,V1679C431,C431V278,C431V611,C431V952,C431V983,C431V1583,C431V1679:std_logic_vector(8 downto 0);
signal V279C432,V612C432,V953C432,V984C432,V1584C432,V1680C432,C432V279,C432V612,C432V953,C432V984,C432V1584,C432V1680:std_logic_vector(8 downto 0);
signal V280C433,V613C433,V954C433,V985C433,V1585C433,V1681C433,C433V280,C433V613,C433V954,C433V985,C433V1585,C433V1681:std_logic_vector(8 downto 0);
signal V281C434,V614C434,V955C434,V986C434,V1586C434,V1682C434,C434V281,C434V614,C434V955,C434V986,C434V1586,C434V1682:std_logic_vector(8 downto 0);
signal V282C435,V615C435,V956C435,V987C435,V1587C435,V1683C435,C435V282,C435V615,C435V956,C435V987,C435V1587,C435V1683:std_logic_vector(8 downto 0);
signal V283C436,V616C436,V957C436,V988C436,V1588C436,V1684C436,C436V283,C436V616,C436V957,C436V988,C436V1588,C436V1684:std_logic_vector(8 downto 0);
signal V284C437,V617C437,V958C437,V989C437,V1589C437,V1685C437,C437V284,C437V617,C437V958,C437V989,C437V1589,C437V1685:std_logic_vector(8 downto 0);
signal V285C438,V618C438,V959C438,V990C438,V1590C438,V1686C438,C438V285,C438V618,C438V959,C438V990,C438V1590,C438V1686:std_logic_vector(8 downto 0);
signal V286C439,V619C439,V960C439,V991C439,V1591C439,V1687C439,C439V286,C439V619,C439V960,C439V991,C439V1591,C439V1687:std_logic_vector(8 downto 0);
signal V287C440,V620C440,V865C440,V992C440,V1592C440,V1688C440,C440V287,C440V620,C440V865,C440V992,C440V1592,C440V1688:std_logic_vector(8 downto 0);
signal V288C441,V621C441,V866C441,V993C441,V1593C441,V1689C441,C441V288,C441V621,C441V866,C441V993,C441V1593,C441V1689:std_logic_vector(8 downto 0);
signal V193C442,V622C442,V867C442,V994C442,V1594C442,V1690C442,C442V193,C442V622,C442V867,C442V994,C442V1594,C442V1690:std_logic_vector(8 downto 0);
signal V194C443,V623C443,V868C443,V995C443,V1595C443,V1691C443,C443V194,C443V623,C443V868,C443V995,C443V1595,C443V1691:std_logic_vector(8 downto 0);
signal V195C444,V624C444,V869C444,V996C444,V1596C444,V1692C444,C444V195,C444V624,C444V869,C444V996,C444V1596,C444V1692:std_logic_vector(8 downto 0);
signal V196C445,V625C445,V870C445,V997C445,V1597C445,V1693C445,C445V196,C445V625,C445V870,C445V997,C445V1597,C445V1693:std_logic_vector(8 downto 0);
signal V197C446,V626C446,V871C446,V998C446,V1598C446,V1694C446,C446V197,C446V626,C446V871,C446V998,C446V1598,C446V1694:std_logic_vector(8 downto 0);
signal V198C447,V627C447,V872C447,V999C447,V1599C447,V1695C447,C447V198,C447V627,C447V872,C447V999,C447V1599,C447V1695:std_logic_vector(8 downto 0);
signal V199C448,V628C448,V873C448,V1000C448,V1600C448,V1696C448,C448V199,C448V628,C448V873,C448V1000,C448V1600,C448V1696:std_logic_vector(8 downto 0);
signal V200C449,V629C449,V874C449,V1001C449,V1601C449,V1697C449,C449V200,C449V629,C449V874,C449V1001,C449V1601,C449V1697:std_logic_vector(8 downto 0);
signal V201C450,V630C450,V875C450,V1002C450,V1602C450,V1698C450,C450V201,C450V630,C450V875,C450V1002,C450V1602,C450V1698:std_logic_vector(8 downto 0);
signal V202C451,V631C451,V876C451,V1003C451,V1603C451,V1699C451,C451V202,C451V631,C451V876,C451V1003,C451V1603,C451V1699:std_logic_vector(8 downto 0);
signal V203C452,V632C452,V877C452,V1004C452,V1604C452,V1700C452,C452V203,C452V632,C452V877,C452V1004,C452V1604,C452V1700:std_logic_vector(8 downto 0);
signal V204C453,V633C453,V878C453,V1005C453,V1605C453,V1701C453,C453V204,C453V633,C453V878,C453V1005,C453V1605,C453V1701:std_logic_vector(8 downto 0);
signal V205C454,V634C454,V879C454,V1006C454,V1606C454,V1702C454,C454V205,C454V634,C454V879,C454V1006,C454V1606,C454V1702:std_logic_vector(8 downto 0);
signal V206C455,V635C455,V880C455,V1007C455,V1607C455,V1703C455,C455V206,C455V635,C455V880,C455V1007,C455V1607,C455V1703:std_logic_vector(8 downto 0);
signal V207C456,V636C456,V881C456,V1008C456,V1608C456,V1704C456,C456V207,C456V636,C456V881,C456V1008,C456V1608,C456V1704:std_logic_vector(8 downto 0);
signal V208C457,V637C457,V882C457,V1009C457,V1609C457,V1705C457,C457V208,C457V637,C457V882,C457V1009,C457V1609,C457V1705:std_logic_vector(8 downto 0);
signal V209C458,V638C458,V883C458,V1010C458,V1610C458,V1706C458,C458V209,C458V638,C458V883,C458V1010,C458V1610,C458V1706:std_logic_vector(8 downto 0);
signal V210C459,V639C459,V884C459,V1011C459,V1611C459,V1707C459,C459V210,C459V639,C459V884,C459V1011,C459V1611,C459V1707:std_logic_vector(8 downto 0);
signal V211C460,V640C460,V885C460,V1012C460,V1612C460,V1708C460,C460V211,C460V640,C460V885,C460V1012,C460V1612,C460V1708:std_logic_vector(8 downto 0);
signal V212C461,V641C461,V886C461,V1013C461,V1613C461,V1709C461,C461V212,C461V641,C461V886,C461V1013,C461V1613,C461V1709:std_logic_vector(8 downto 0);
signal V213C462,V642C462,V887C462,V1014C462,V1614C462,V1710C462,C462V213,C462V642,C462V887,C462V1014,C462V1614,C462V1710:std_logic_vector(8 downto 0);
signal V214C463,V643C463,V888C463,V1015C463,V1615C463,V1711C463,C463V214,C463V643,C463V888,C463V1015,C463V1615,C463V1711:std_logic_vector(8 downto 0);
signal V215C464,V644C464,V889C464,V1016C464,V1616C464,V1712C464,C464V215,C464V644,C464V889,C464V1016,C464V1616,C464V1712:std_logic_vector(8 downto 0);
signal V216C465,V645C465,V890C465,V1017C465,V1617C465,V1713C465,C465V216,C465V645,C465V890,C465V1017,C465V1617,C465V1713:std_logic_vector(8 downto 0);
signal V217C466,V646C466,V891C466,V1018C466,V1618C466,V1714C466,C466V217,C466V646,C466V891,C466V1018,C466V1618,C466V1714:std_logic_vector(8 downto 0);
signal V218C467,V647C467,V892C467,V1019C467,V1619C467,V1715C467,C467V218,C467V647,C467V892,C467V1019,C467V1619,C467V1715:std_logic_vector(8 downto 0);
signal V219C468,V648C468,V893C468,V1020C468,V1620C468,V1716C468,C468V219,C468V648,C468V893,C468V1020,C468V1620,C468V1716:std_logic_vector(8 downto 0);
signal V220C469,V649C469,V894C469,V1021C469,V1621C469,V1717C469,C469V220,C469V649,C469V894,C469V1021,C469V1621,C469V1717:std_logic_vector(8 downto 0);
signal V221C470,V650C470,V895C470,V1022C470,V1622C470,V1718C470,C470V221,C470V650,C470V895,C470V1022,C470V1622,C470V1718:std_logic_vector(8 downto 0);
signal V222C471,V651C471,V896C471,V1023C471,V1623C471,V1719C471,C471V222,C471V651,C471V896,C471V1023,C471V1623,C471V1719:std_logic_vector(8 downto 0);
signal V223C472,V652C472,V897C472,V1024C472,V1624C472,V1720C472,C472V223,C472V652,C472V897,C472V1024,C472V1624,C472V1720:std_logic_vector(8 downto 0);
signal V224C473,V653C473,V898C473,V1025C473,V1625C473,V1721C473,C473V224,C473V653,C473V898,C473V1025,C473V1625,C473V1721:std_logic_vector(8 downto 0);
signal V225C474,V654C474,V899C474,V1026C474,V1626C474,V1722C474,C474V225,C474V654,C474V899,C474V1026,C474V1626,C474V1722:std_logic_vector(8 downto 0);
signal V226C475,V655C475,V900C475,V1027C475,V1627C475,V1723C475,C475V226,C475V655,C475V900,C475V1027,C475V1627,C475V1723:std_logic_vector(8 downto 0);
signal V227C476,V656C476,V901C476,V1028C476,V1628C476,V1724C476,C476V227,C476V656,C476V901,C476V1028,C476V1628,C476V1724:std_logic_vector(8 downto 0);
signal V228C477,V657C477,V902C477,V1029C477,V1629C477,V1725C477,C477V228,C477V657,C477V902,C477V1029,C477V1629,C477V1725:std_logic_vector(8 downto 0);
signal V229C478,V658C478,V903C478,V1030C478,V1630C478,V1726C478,C478V229,C478V658,C478V903,C478V1030,C478V1630,C478V1726:std_logic_vector(8 downto 0);
signal V230C479,V659C479,V904C479,V1031C479,V1631C479,V1727C479,C479V230,C479V659,C479V904,C479V1031,C479V1631,C479V1727:std_logic_vector(8 downto 0);
signal V231C480,V660C480,V905C480,V1032C480,V1632C480,V1728C480,C480V231,C480V660,C480V905,C480V1032,C480V1632,C480V1728:std_logic_vector(8 downto 0);
signal V431C481,V521C481,V755C481,V1136C481,V1153C481,V1633C481,V1729C481,C481V431,C481V521,C481V755,C481V1136,C481V1153,C481V1633,C481V1729:std_logic_vector(8 downto 0);
signal V432C482,V522C482,V756C482,V1137C482,V1154C482,V1634C482,V1730C482,C482V432,C482V522,C482V756,C482V1137,C482V1154,C482V1634,C482V1730:std_logic_vector(8 downto 0);
signal V433C483,V523C483,V757C483,V1138C483,V1155C483,V1635C483,V1731C483,C483V433,C483V523,C483V757,C483V1138,C483V1155,C483V1635,C483V1731:std_logic_vector(8 downto 0);
signal V434C484,V524C484,V758C484,V1139C484,V1156C484,V1636C484,V1732C484,C484V434,C484V524,C484V758,C484V1139,C484V1156,C484V1636,C484V1732:std_logic_vector(8 downto 0);
signal V435C485,V525C485,V759C485,V1140C485,V1157C485,V1637C485,V1733C485,C485V435,C485V525,C485V759,C485V1140,C485V1157,C485V1637,C485V1733:std_logic_vector(8 downto 0);
signal V436C486,V526C486,V760C486,V1141C486,V1158C486,V1638C486,V1734C486,C486V436,C486V526,C486V760,C486V1141,C486V1158,C486V1638,C486V1734:std_logic_vector(8 downto 0);
signal V437C487,V527C487,V761C487,V1142C487,V1159C487,V1639C487,V1735C487,C487V437,C487V527,C487V761,C487V1142,C487V1159,C487V1639,C487V1735:std_logic_vector(8 downto 0);
signal V438C488,V528C488,V762C488,V1143C488,V1160C488,V1640C488,V1736C488,C488V438,C488V528,C488V762,C488V1143,C488V1160,C488V1640,C488V1736:std_logic_vector(8 downto 0);
signal V439C489,V529C489,V763C489,V1144C489,V1161C489,V1641C489,V1737C489,C489V439,C489V529,C489V763,C489V1144,C489V1161,C489V1641,C489V1737:std_logic_vector(8 downto 0);
signal V440C490,V530C490,V764C490,V1145C490,V1162C490,V1642C490,V1738C490,C490V440,C490V530,C490V764,C490V1145,C490V1162,C490V1642,C490V1738:std_logic_vector(8 downto 0);
signal V441C491,V531C491,V765C491,V1146C491,V1163C491,V1643C491,V1739C491,C491V441,C491V531,C491V765,C491V1146,C491V1163,C491V1643,C491V1739:std_logic_vector(8 downto 0);
signal V442C492,V532C492,V766C492,V1147C492,V1164C492,V1644C492,V1740C492,C492V442,C492V532,C492V766,C492V1147,C492V1164,C492V1644,C492V1740:std_logic_vector(8 downto 0);
signal V443C493,V533C493,V767C493,V1148C493,V1165C493,V1645C493,V1741C493,C493V443,C493V533,C493V767,C493V1148,C493V1165,C493V1645,C493V1741:std_logic_vector(8 downto 0);
signal V444C494,V534C494,V768C494,V1149C494,V1166C494,V1646C494,V1742C494,C494V444,C494V534,C494V768,C494V1149,C494V1166,C494V1646,C494V1742:std_logic_vector(8 downto 0);
signal V445C495,V535C495,V673C495,V1150C495,V1167C495,V1647C495,V1743C495,C495V445,C495V535,C495V673,C495V1150,C495V1167,C495V1647,C495V1743:std_logic_vector(8 downto 0);
signal V446C496,V536C496,V674C496,V1151C496,V1168C496,V1648C496,V1744C496,C496V446,C496V536,C496V674,C496V1151,C496V1168,C496V1648,C496V1744:std_logic_vector(8 downto 0);
signal V447C497,V537C497,V675C497,V1152C497,V1169C497,V1649C497,V1745C497,C497V447,C497V537,C497V675,C497V1152,C497V1169,C497V1649,C497V1745:std_logic_vector(8 downto 0);
signal V448C498,V538C498,V676C498,V1057C498,V1170C498,V1650C498,V1746C498,C498V448,C498V538,C498V676,C498V1057,C498V1170,C498V1650,C498V1746:std_logic_vector(8 downto 0);
signal V449C499,V539C499,V677C499,V1058C499,V1171C499,V1651C499,V1747C499,C499V449,C499V539,C499V677,C499V1058,C499V1171,C499V1651,C499V1747:std_logic_vector(8 downto 0);
signal V450C500,V540C500,V678C500,V1059C500,V1172C500,V1652C500,V1748C500,C500V450,C500V540,C500V678,C500V1059,C500V1172,C500V1652,C500V1748:std_logic_vector(8 downto 0);
signal V451C501,V541C501,V679C501,V1060C501,V1173C501,V1653C501,V1749C501,C501V451,C501V541,C501V679,C501V1060,C501V1173,C501V1653,C501V1749:std_logic_vector(8 downto 0);
signal V452C502,V542C502,V680C502,V1061C502,V1174C502,V1654C502,V1750C502,C502V452,C502V542,C502V680,C502V1061,C502V1174,C502V1654,C502V1750:std_logic_vector(8 downto 0);
signal V453C503,V543C503,V681C503,V1062C503,V1175C503,V1655C503,V1751C503,C503V453,C503V543,C503V681,C503V1062,C503V1175,C503V1655,C503V1751:std_logic_vector(8 downto 0);
signal V454C504,V544C504,V682C504,V1063C504,V1176C504,V1656C504,V1752C504,C504V454,C504V544,C504V682,C504V1063,C504V1176,C504V1656,C504V1752:std_logic_vector(8 downto 0);
signal V455C505,V545C505,V683C505,V1064C505,V1177C505,V1657C505,V1753C505,C505V455,C505V545,C505V683,C505V1064,C505V1177,C505V1657,C505V1753:std_logic_vector(8 downto 0);
signal V456C506,V546C506,V684C506,V1065C506,V1178C506,V1658C506,V1754C506,C506V456,C506V546,C506V684,C506V1065,C506V1178,C506V1658,C506V1754:std_logic_vector(8 downto 0);
signal V457C507,V547C507,V685C507,V1066C507,V1179C507,V1659C507,V1755C507,C507V457,C507V547,C507V685,C507V1066,C507V1179,C507V1659,C507V1755:std_logic_vector(8 downto 0);
signal V458C508,V548C508,V686C508,V1067C508,V1180C508,V1660C508,V1756C508,C508V458,C508V548,C508V686,C508V1067,C508V1180,C508V1660,C508V1756:std_logic_vector(8 downto 0);
signal V459C509,V549C509,V687C509,V1068C509,V1181C509,V1661C509,V1757C509,C509V459,C509V549,C509V687,C509V1068,C509V1181,C509V1661,C509V1757:std_logic_vector(8 downto 0);
signal V460C510,V550C510,V688C510,V1069C510,V1182C510,V1662C510,V1758C510,C510V460,C510V550,C510V688,C510V1069,C510V1182,C510V1662,C510V1758:std_logic_vector(8 downto 0);
signal V461C511,V551C511,V689C511,V1070C511,V1183C511,V1663C511,V1759C511,C511V461,C511V551,C511V689,C511V1070,C511V1183,C511V1663,C511V1759:std_logic_vector(8 downto 0);
signal V462C512,V552C512,V690C512,V1071C512,V1184C512,V1664C512,V1760C512,C512V462,C512V552,C512V690,C512V1071,C512V1184,C512V1664,C512V1760:std_logic_vector(8 downto 0);
signal V463C513,V553C513,V691C513,V1072C513,V1185C513,V1665C513,V1761C513,C513V463,C513V553,C513V691,C513V1072,C513V1185,C513V1665,C513V1761:std_logic_vector(8 downto 0);
signal V464C514,V554C514,V692C514,V1073C514,V1186C514,V1666C514,V1762C514,C514V464,C514V554,C514V692,C514V1073,C514V1186,C514V1666,C514V1762:std_logic_vector(8 downto 0);
signal V465C515,V555C515,V693C515,V1074C515,V1187C515,V1667C515,V1763C515,C515V465,C515V555,C515V693,C515V1074,C515V1187,C515V1667,C515V1763:std_logic_vector(8 downto 0);
signal V466C516,V556C516,V694C516,V1075C516,V1188C516,V1668C516,V1764C516,C516V466,C516V556,C516V694,C516V1075,C516V1188,C516V1668,C516V1764:std_logic_vector(8 downto 0);
signal V467C517,V557C517,V695C517,V1076C517,V1189C517,V1669C517,V1765C517,C517V467,C517V557,C517V695,C517V1076,C517V1189,C517V1669,C517V1765:std_logic_vector(8 downto 0);
signal V468C518,V558C518,V696C518,V1077C518,V1190C518,V1670C518,V1766C518,C518V468,C518V558,C518V696,C518V1077,C518V1190,C518V1670,C518V1766:std_logic_vector(8 downto 0);
signal V469C519,V559C519,V697C519,V1078C519,V1191C519,V1671C519,V1767C519,C519V469,C519V559,C519V697,C519V1078,C519V1191,C519V1671,C519V1767:std_logic_vector(8 downto 0);
signal V470C520,V560C520,V698C520,V1079C520,V1192C520,V1672C520,V1768C520,C520V470,C520V560,C520V698,C520V1079,C520V1192,C520V1672,C520V1768:std_logic_vector(8 downto 0);
signal V471C521,V561C521,V699C521,V1080C521,V1193C521,V1673C521,V1769C521,C521V471,C521V561,C521V699,C521V1080,C521V1193,C521V1673,C521V1769:std_logic_vector(8 downto 0);
signal V472C522,V562C522,V700C522,V1081C522,V1194C522,V1674C522,V1770C522,C522V472,C522V562,C522V700,C522V1081,C522V1194,C522V1674,C522V1770:std_logic_vector(8 downto 0);
signal V473C523,V563C523,V701C523,V1082C523,V1195C523,V1675C523,V1771C523,C523V473,C523V563,C523V701,C523V1082,C523V1195,C523V1675,C523V1771:std_logic_vector(8 downto 0);
signal V474C524,V564C524,V702C524,V1083C524,V1196C524,V1676C524,V1772C524,C524V474,C524V564,C524V702,C524V1083,C524V1196,C524V1676,C524V1772:std_logic_vector(8 downto 0);
signal V475C525,V565C525,V703C525,V1084C525,V1197C525,V1677C525,V1773C525,C525V475,C525V565,C525V703,C525V1084,C525V1197,C525V1677,C525V1773:std_logic_vector(8 downto 0);
signal V476C526,V566C526,V704C526,V1085C526,V1198C526,V1678C526,V1774C526,C526V476,C526V566,C526V704,C526V1085,C526V1198,C526V1678,C526V1774:std_logic_vector(8 downto 0);
signal V477C527,V567C527,V705C527,V1086C527,V1199C527,V1679C527,V1775C527,C527V477,C527V567,C527V705,C527V1086,C527V1199,C527V1679,C527V1775:std_logic_vector(8 downto 0);
signal V478C528,V568C528,V706C528,V1087C528,V1200C528,V1680C528,V1776C528,C528V478,C528V568,C528V706,C528V1087,C528V1200,C528V1680,C528V1776:std_logic_vector(8 downto 0);
signal V479C529,V569C529,V707C529,V1088C529,V1201C529,V1681C529,V1777C529,C529V479,C529V569,C529V707,C529V1088,C529V1201,C529V1681,C529V1777:std_logic_vector(8 downto 0);
signal V480C530,V570C530,V708C530,V1089C530,V1202C530,V1682C530,V1778C530,C530V480,C530V570,C530V708,C530V1089,C530V1202,C530V1682,C530V1778:std_logic_vector(8 downto 0);
signal V385C531,V571C531,V709C531,V1090C531,V1203C531,V1683C531,V1779C531,C531V385,C531V571,C531V709,C531V1090,C531V1203,C531V1683,C531V1779:std_logic_vector(8 downto 0);
signal V386C532,V572C532,V710C532,V1091C532,V1204C532,V1684C532,V1780C532,C532V386,C532V572,C532V710,C532V1091,C532V1204,C532V1684,C532V1780:std_logic_vector(8 downto 0);
signal V387C533,V573C533,V711C533,V1092C533,V1205C533,V1685C533,V1781C533,C533V387,C533V573,C533V711,C533V1092,C533V1205,C533V1685,C533V1781:std_logic_vector(8 downto 0);
signal V388C534,V574C534,V712C534,V1093C534,V1206C534,V1686C534,V1782C534,C534V388,C534V574,C534V712,C534V1093,C534V1206,C534V1686,C534V1782:std_logic_vector(8 downto 0);
signal V389C535,V575C535,V713C535,V1094C535,V1207C535,V1687C535,V1783C535,C535V389,C535V575,C535V713,C535V1094,C535V1207,C535V1687,C535V1783:std_logic_vector(8 downto 0);
signal V390C536,V576C536,V714C536,V1095C536,V1208C536,V1688C536,V1784C536,C536V390,C536V576,C536V714,C536V1095,C536V1208,C536V1688,C536V1784:std_logic_vector(8 downto 0);
signal V391C537,V481C537,V715C537,V1096C537,V1209C537,V1689C537,V1785C537,C537V391,C537V481,C537V715,C537V1096,C537V1209,C537V1689,C537V1785:std_logic_vector(8 downto 0);
signal V392C538,V482C538,V716C538,V1097C538,V1210C538,V1690C538,V1786C538,C538V392,C538V482,C538V716,C538V1097,C538V1210,C538V1690,C538V1786:std_logic_vector(8 downto 0);
signal V393C539,V483C539,V717C539,V1098C539,V1211C539,V1691C539,V1787C539,C539V393,C539V483,C539V717,C539V1098,C539V1211,C539V1691,C539V1787:std_logic_vector(8 downto 0);
signal V394C540,V484C540,V718C540,V1099C540,V1212C540,V1692C540,V1788C540,C540V394,C540V484,C540V718,C540V1099,C540V1212,C540V1692,C540V1788:std_logic_vector(8 downto 0);
signal V395C541,V485C541,V719C541,V1100C541,V1213C541,V1693C541,V1789C541,C541V395,C541V485,C541V719,C541V1100,C541V1213,C541V1693,C541V1789:std_logic_vector(8 downto 0);
signal V396C542,V486C542,V720C542,V1101C542,V1214C542,V1694C542,V1790C542,C542V396,C542V486,C542V720,C542V1101,C542V1214,C542V1694,C542V1790:std_logic_vector(8 downto 0);
signal V397C543,V487C543,V721C543,V1102C543,V1215C543,V1695C543,V1791C543,C543V397,C543V487,C543V721,C543V1102,C543V1215,C543V1695,C543V1791:std_logic_vector(8 downto 0);
signal V398C544,V488C544,V722C544,V1103C544,V1216C544,V1696C544,V1792C544,C544V398,C544V488,C544V722,C544V1103,C544V1216,C544V1696,C544V1792:std_logic_vector(8 downto 0);
signal V399C545,V489C545,V723C545,V1104C545,V1217C545,V1697C545,V1793C545,C545V399,C545V489,C545V723,C545V1104,C545V1217,C545V1697,C545V1793:std_logic_vector(8 downto 0);
signal V400C546,V490C546,V724C546,V1105C546,V1218C546,V1698C546,V1794C546,C546V400,C546V490,C546V724,C546V1105,C546V1218,C546V1698,C546V1794:std_logic_vector(8 downto 0);
signal V401C547,V491C547,V725C547,V1106C547,V1219C547,V1699C547,V1795C547,C547V401,C547V491,C547V725,C547V1106,C547V1219,C547V1699,C547V1795:std_logic_vector(8 downto 0);
signal V402C548,V492C548,V726C548,V1107C548,V1220C548,V1700C548,V1796C548,C548V402,C548V492,C548V726,C548V1107,C548V1220,C548V1700,C548V1796:std_logic_vector(8 downto 0);
signal V403C549,V493C549,V727C549,V1108C549,V1221C549,V1701C549,V1797C549,C549V403,C549V493,C549V727,C549V1108,C549V1221,C549V1701,C549V1797:std_logic_vector(8 downto 0);
signal V404C550,V494C550,V728C550,V1109C550,V1222C550,V1702C550,V1798C550,C550V404,C550V494,C550V728,C550V1109,C550V1222,C550V1702,C550V1798:std_logic_vector(8 downto 0);
signal V405C551,V495C551,V729C551,V1110C551,V1223C551,V1703C551,V1799C551,C551V405,C551V495,C551V729,C551V1110,C551V1223,C551V1703,C551V1799:std_logic_vector(8 downto 0);
signal V406C552,V496C552,V730C552,V1111C552,V1224C552,V1704C552,V1800C552,C552V406,C552V496,C552V730,C552V1111,C552V1224,C552V1704,C552V1800:std_logic_vector(8 downto 0);
signal V407C553,V497C553,V731C553,V1112C553,V1225C553,V1705C553,V1801C553,C553V407,C553V497,C553V731,C553V1112,C553V1225,C553V1705,C553V1801:std_logic_vector(8 downto 0);
signal V408C554,V498C554,V732C554,V1113C554,V1226C554,V1706C554,V1802C554,C554V408,C554V498,C554V732,C554V1113,C554V1226,C554V1706,C554V1802:std_logic_vector(8 downto 0);
signal V409C555,V499C555,V733C555,V1114C555,V1227C555,V1707C555,V1803C555,C555V409,C555V499,C555V733,C555V1114,C555V1227,C555V1707,C555V1803:std_logic_vector(8 downto 0);
signal V410C556,V500C556,V734C556,V1115C556,V1228C556,V1708C556,V1804C556,C556V410,C556V500,C556V734,C556V1115,C556V1228,C556V1708,C556V1804:std_logic_vector(8 downto 0);
signal V411C557,V501C557,V735C557,V1116C557,V1229C557,V1709C557,V1805C557,C557V411,C557V501,C557V735,C557V1116,C557V1229,C557V1709,C557V1805:std_logic_vector(8 downto 0);
signal V412C558,V502C558,V736C558,V1117C558,V1230C558,V1710C558,V1806C558,C558V412,C558V502,C558V736,C558V1117,C558V1230,C558V1710,C558V1806:std_logic_vector(8 downto 0);
signal V413C559,V503C559,V737C559,V1118C559,V1231C559,V1711C559,V1807C559,C559V413,C559V503,C559V737,C559V1118,C559V1231,C559V1711,C559V1807:std_logic_vector(8 downto 0);
signal V414C560,V504C560,V738C560,V1119C560,V1232C560,V1712C560,V1808C560,C560V414,C560V504,C560V738,C560V1119,C560V1232,C560V1712,C560V1808:std_logic_vector(8 downto 0);
signal V415C561,V505C561,V739C561,V1120C561,V1233C561,V1713C561,V1809C561,C561V415,C561V505,C561V739,C561V1120,C561V1233,C561V1713,C561V1809:std_logic_vector(8 downto 0);
signal V416C562,V506C562,V740C562,V1121C562,V1234C562,V1714C562,V1810C562,C562V416,C562V506,C562V740,C562V1121,C562V1234,C562V1714,C562V1810:std_logic_vector(8 downto 0);
signal V417C563,V507C563,V741C563,V1122C563,V1235C563,V1715C563,V1811C563,C563V417,C563V507,C563V741,C563V1122,C563V1235,C563V1715,C563V1811:std_logic_vector(8 downto 0);
signal V418C564,V508C564,V742C564,V1123C564,V1236C564,V1716C564,V1812C564,C564V418,C564V508,C564V742,C564V1123,C564V1236,C564V1716,C564V1812:std_logic_vector(8 downto 0);
signal V419C565,V509C565,V743C565,V1124C565,V1237C565,V1717C565,V1813C565,C565V419,C565V509,C565V743,C565V1124,C565V1237,C565V1717,C565V1813:std_logic_vector(8 downto 0);
signal V420C566,V510C566,V744C566,V1125C566,V1238C566,V1718C566,V1814C566,C566V420,C566V510,C566V744,C566V1125,C566V1238,C566V1718,C566V1814:std_logic_vector(8 downto 0);
signal V421C567,V511C567,V745C567,V1126C567,V1239C567,V1719C567,V1815C567,C567V421,C567V511,C567V745,C567V1126,C567V1239,C567V1719,C567V1815:std_logic_vector(8 downto 0);
signal V422C568,V512C568,V746C568,V1127C568,V1240C568,V1720C568,V1816C568,C568V422,C568V512,C568V746,C568V1127,C568V1240,C568V1720,C568V1816:std_logic_vector(8 downto 0);
signal V423C569,V513C569,V747C569,V1128C569,V1241C569,V1721C569,V1817C569,C569V423,C569V513,C569V747,C569V1128,C569V1241,C569V1721,C569V1817:std_logic_vector(8 downto 0);
signal V424C570,V514C570,V748C570,V1129C570,V1242C570,V1722C570,V1818C570,C570V424,C570V514,C570V748,C570V1129,C570V1242,C570V1722,C570V1818:std_logic_vector(8 downto 0);
signal V425C571,V515C571,V749C571,V1130C571,V1243C571,V1723C571,V1819C571,C571V425,C571V515,C571V749,C571V1130,C571V1243,C571V1723,C571V1819:std_logic_vector(8 downto 0);
signal V426C572,V516C572,V750C572,V1131C572,V1244C572,V1724C572,V1820C572,C572V426,C572V516,C572V750,C572V1131,C572V1244,C572V1724,C572V1820:std_logic_vector(8 downto 0);
signal V427C573,V517C573,V751C573,V1132C573,V1245C573,V1725C573,V1821C573,C573V427,C573V517,C573V751,C573V1132,C573V1245,C573V1725,C573V1821:std_logic_vector(8 downto 0);
signal V428C574,V518C574,V752C574,V1133C574,V1246C574,V1726C574,V1822C574,C574V428,C574V518,C574V752,C574V1133,C574V1246,C574V1726,C574V1822:std_logic_vector(8 downto 0);
signal V429C575,V519C575,V753C575,V1134C575,V1247C575,V1727C575,V1823C575,C575V429,C575V519,C575V753,C575V1134,C575V1247,C575V1727,C575V1823:std_logic_vector(8 downto 0);
signal V430C576,V520C576,V754C576,V1135C576,V1248C576,V1728C576,V1824C576,C576V430,C576V520,C576V754,C576V1135,C576V1248,C576V1728,C576V1824:std_logic_vector(8 downto 0);
signal V288C577,V342C577,V879C577,V979C577,V1729C577,V1825C577,C577V288,C577V342,C577V879,C577V979,C577V1729,C577V1825:std_logic_vector(8 downto 0);
signal V193C578,V343C578,V880C578,V980C578,V1730C578,V1826C578,C578V193,C578V343,C578V880,C578V980,C578V1730,C578V1826:std_logic_vector(8 downto 0);
signal V194C579,V344C579,V881C579,V981C579,V1731C579,V1827C579,C579V194,C579V344,C579V881,C579V981,C579V1731,C579V1827:std_logic_vector(8 downto 0);
signal V195C580,V345C580,V882C580,V982C580,V1732C580,V1828C580,C580V195,C580V345,C580V882,C580V982,C580V1732,C580V1828:std_logic_vector(8 downto 0);
signal V196C581,V346C581,V883C581,V983C581,V1733C581,V1829C581,C581V196,C581V346,C581V883,C581V983,C581V1733,C581V1829:std_logic_vector(8 downto 0);
signal V197C582,V347C582,V884C582,V984C582,V1734C582,V1830C582,C582V197,C582V347,C582V884,C582V984,C582V1734,C582V1830:std_logic_vector(8 downto 0);
signal V198C583,V348C583,V885C583,V985C583,V1735C583,V1831C583,C583V198,C583V348,C583V885,C583V985,C583V1735,C583V1831:std_logic_vector(8 downto 0);
signal V199C584,V349C584,V886C584,V986C584,V1736C584,V1832C584,C584V199,C584V349,C584V886,C584V986,C584V1736,C584V1832:std_logic_vector(8 downto 0);
signal V200C585,V350C585,V887C585,V987C585,V1737C585,V1833C585,C585V200,C585V350,C585V887,C585V987,C585V1737,C585V1833:std_logic_vector(8 downto 0);
signal V201C586,V351C586,V888C586,V988C586,V1738C586,V1834C586,C586V201,C586V351,C586V888,C586V988,C586V1738,C586V1834:std_logic_vector(8 downto 0);
signal V202C587,V352C587,V889C587,V989C587,V1739C587,V1835C587,C587V202,C587V352,C587V889,C587V989,C587V1739,C587V1835:std_logic_vector(8 downto 0);
signal V203C588,V353C588,V890C588,V990C588,V1740C588,V1836C588,C588V203,C588V353,C588V890,C588V990,C588V1740,C588V1836:std_logic_vector(8 downto 0);
signal V204C589,V354C589,V891C589,V991C589,V1741C589,V1837C589,C589V204,C589V354,C589V891,C589V991,C589V1741,C589V1837:std_logic_vector(8 downto 0);
signal V205C590,V355C590,V892C590,V992C590,V1742C590,V1838C590,C590V205,C590V355,C590V892,C590V992,C590V1742,C590V1838:std_logic_vector(8 downto 0);
signal V206C591,V356C591,V893C591,V993C591,V1743C591,V1839C591,C591V206,C591V356,C591V893,C591V993,C591V1743,C591V1839:std_logic_vector(8 downto 0);
signal V207C592,V357C592,V894C592,V994C592,V1744C592,V1840C592,C592V207,C592V357,C592V894,C592V994,C592V1744,C592V1840:std_logic_vector(8 downto 0);
signal V208C593,V358C593,V895C593,V995C593,V1745C593,V1841C593,C593V208,C593V358,C593V895,C593V995,C593V1745,C593V1841:std_logic_vector(8 downto 0);
signal V209C594,V359C594,V896C594,V996C594,V1746C594,V1842C594,C594V209,C594V359,C594V896,C594V996,C594V1746,C594V1842:std_logic_vector(8 downto 0);
signal V210C595,V360C595,V897C595,V997C595,V1747C595,V1843C595,C595V210,C595V360,C595V897,C595V997,C595V1747,C595V1843:std_logic_vector(8 downto 0);
signal V211C596,V361C596,V898C596,V998C596,V1748C596,V1844C596,C596V211,C596V361,C596V898,C596V998,C596V1748,C596V1844:std_logic_vector(8 downto 0);
signal V212C597,V362C597,V899C597,V999C597,V1749C597,V1845C597,C597V212,C597V362,C597V899,C597V999,C597V1749,C597V1845:std_logic_vector(8 downto 0);
signal V213C598,V363C598,V900C598,V1000C598,V1750C598,V1846C598,C598V213,C598V363,C598V900,C598V1000,C598V1750,C598V1846:std_logic_vector(8 downto 0);
signal V214C599,V364C599,V901C599,V1001C599,V1751C599,V1847C599,C599V214,C599V364,C599V901,C599V1001,C599V1751,C599V1847:std_logic_vector(8 downto 0);
signal V215C600,V365C600,V902C600,V1002C600,V1752C600,V1848C600,C600V215,C600V365,C600V902,C600V1002,C600V1752,C600V1848:std_logic_vector(8 downto 0);
signal V216C601,V366C601,V903C601,V1003C601,V1753C601,V1849C601,C601V216,C601V366,C601V903,C601V1003,C601V1753,C601V1849:std_logic_vector(8 downto 0);
signal V217C602,V367C602,V904C602,V1004C602,V1754C602,V1850C602,C602V217,C602V367,C602V904,C602V1004,C602V1754,C602V1850:std_logic_vector(8 downto 0);
signal V218C603,V368C603,V905C603,V1005C603,V1755C603,V1851C603,C603V218,C603V368,C603V905,C603V1005,C603V1755,C603V1851:std_logic_vector(8 downto 0);
signal V219C604,V369C604,V906C604,V1006C604,V1756C604,V1852C604,C604V219,C604V369,C604V906,C604V1006,C604V1756,C604V1852:std_logic_vector(8 downto 0);
signal V220C605,V370C605,V907C605,V1007C605,V1757C605,V1853C605,C605V220,C605V370,C605V907,C605V1007,C605V1757,C605V1853:std_logic_vector(8 downto 0);
signal V221C606,V371C606,V908C606,V1008C606,V1758C606,V1854C606,C606V221,C606V371,C606V908,C606V1008,C606V1758,C606V1854:std_logic_vector(8 downto 0);
signal V222C607,V372C607,V909C607,V1009C607,V1759C607,V1855C607,C607V222,C607V372,C607V909,C607V1009,C607V1759,C607V1855:std_logic_vector(8 downto 0);
signal V223C608,V373C608,V910C608,V1010C608,V1760C608,V1856C608,C608V223,C608V373,C608V910,C608V1010,C608V1760,C608V1856:std_logic_vector(8 downto 0);
signal V224C609,V374C609,V911C609,V1011C609,V1761C609,V1857C609,C609V224,C609V374,C609V911,C609V1011,C609V1761,C609V1857:std_logic_vector(8 downto 0);
signal V225C610,V375C610,V912C610,V1012C610,V1762C610,V1858C610,C610V225,C610V375,C610V912,C610V1012,C610V1762,C610V1858:std_logic_vector(8 downto 0);
signal V226C611,V376C611,V913C611,V1013C611,V1763C611,V1859C611,C611V226,C611V376,C611V913,C611V1013,C611V1763,C611V1859:std_logic_vector(8 downto 0);
signal V227C612,V377C612,V914C612,V1014C612,V1764C612,V1860C612,C612V227,C612V377,C612V914,C612V1014,C612V1764,C612V1860:std_logic_vector(8 downto 0);
signal V228C613,V378C613,V915C613,V1015C613,V1765C613,V1861C613,C613V228,C613V378,C613V915,C613V1015,C613V1765,C613V1861:std_logic_vector(8 downto 0);
signal V229C614,V379C614,V916C614,V1016C614,V1766C614,V1862C614,C614V229,C614V379,C614V916,C614V1016,C614V1766,C614V1862:std_logic_vector(8 downto 0);
signal V230C615,V380C615,V917C615,V1017C615,V1767C615,V1863C615,C615V230,C615V380,C615V917,C615V1017,C615V1767,C615V1863:std_logic_vector(8 downto 0);
signal V231C616,V381C616,V918C616,V1018C616,V1768C616,V1864C616,C616V231,C616V381,C616V918,C616V1018,C616V1768,C616V1864:std_logic_vector(8 downto 0);
signal V232C617,V382C617,V919C617,V1019C617,V1769C617,V1865C617,C617V232,C617V382,C617V919,C617V1019,C617V1769,C617V1865:std_logic_vector(8 downto 0);
signal V233C618,V383C618,V920C618,V1020C618,V1770C618,V1866C618,C618V233,C618V383,C618V920,C618V1020,C618V1770,C618V1866:std_logic_vector(8 downto 0);
signal V234C619,V384C619,V921C619,V1021C619,V1771C619,V1867C619,C619V234,C619V384,C619V921,C619V1021,C619V1771,C619V1867:std_logic_vector(8 downto 0);
signal V235C620,V289C620,V922C620,V1022C620,V1772C620,V1868C620,C620V235,C620V289,C620V922,C620V1022,C620V1772,C620V1868:std_logic_vector(8 downto 0);
signal V236C621,V290C621,V923C621,V1023C621,V1773C621,V1869C621,C621V236,C621V290,C621V923,C621V1023,C621V1773,C621V1869:std_logic_vector(8 downto 0);
signal V237C622,V291C622,V924C622,V1024C622,V1774C622,V1870C622,C622V237,C622V291,C622V924,C622V1024,C622V1774,C622V1870:std_logic_vector(8 downto 0);
signal V238C623,V292C623,V925C623,V1025C623,V1775C623,V1871C623,C623V238,C623V292,C623V925,C623V1025,C623V1775,C623V1871:std_logic_vector(8 downto 0);
signal V239C624,V293C624,V926C624,V1026C624,V1776C624,V1872C624,C624V239,C624V293,C624V926,C624V1026,C624V1776,C624V1872:std_logic_vector(8 downto 0);
signal V240C625,V294C625,V927C625,V1027C625,V1777C625,V1873C625,C625V240,C625V294,C625V927,C625V1027,C625V1777,C625V1873:std_logic_vector(8 downto 0);
signal V241C626,V295C626,V928C626,V1028C626,V1778C626,V1874C626,C626V241,C626V295,C626V928,C626V1028,C626V1778,C626V1874:std_logic_vector(8 downto 0);
signal V242C627,V296C627,V929C627,V1029C627,V1779C627,V1875C627,C627V242,C627V296,C627V929,C627V1029,C627V1779,C627V1875:std_logic_vector(8 downto 0);
signal V243C628,V297C628,V930C628,V1030C628,V1780C628,V1876C628,C628V243,C628V297,C628V930,C628V1030,C628V1780,C628V1876:std_logic_vector(8 downto 0);
signal V244C629,V298C629,V931C629,V1031C629,V1781C629,V1877C629,C629V244,C629V298,C629V931,C629V1031,C629V1781,C629V1877:std_logic_vector(8 downto 0);
signal V245C630,V299C630,V932C630,V1032C630,V1782C630,V1878C630,C630V245,C630V299,C630V932,C630V1032,C630V1782,C630V1878:std_logic_vector(8 downto 0);
signal V246C631,V300C631,V933C631,V1033C631,V1783C631,V1879C631,C631V246,C631V300,C631V933,C631V1033,C631V1783,C631V1879:std_logic_vector(8 downto 0);
signal V247C632,V301C632,V934C632,V1034C632,V1784C632,V1880C632,C632V247,C632V301,C632V934,C632V1034,C632V1784,C632V1880:std_logic_vector(8 downto 0);
signal V248C633,V302C633,V935C633,V1035C633,V1785C633,V1881C633,C633V248,C633V302,C633V935,C633V1035,C633V1785,C633V1881:std_logic_vector(8 downto 0);
signal V249C634,V303C634,V936C634,V1036C634,V1786C634,V1882C634,C634V249,C634V303,C634V936,C634V1036,C634V1786,C634V1882:std_logic_vector(8 downto 0);
signal V250C635,V304C635,V937C635,V1037C635,V1787C635,V1883C635,C635V250,C635V304,C635V937,C635V1037,C635V1787,C635V1883:std_logic_vector(8 downto 0);
signal V251C636,V305C636,V938C636,V1038C636,V1788C636,V1884C636,C636V251,C636V305,C636V938,C636V1038,C636V1788,C636V1884:std_logic_vector(8 downto 0);
signal V252C637,V306C637,V939C637,V1039C637,V1789C637,V1885C637,C637V252,C637V306,C637V939,C637V1039,C637V1789,C637V1885:std_logic_vector(8 downto 0);
signal V253C638,V307C638,V940C638,V1040C638,V1790C638,V1886C638,C638V253,C638V307,C638V940,C638V1040,C638V1790,C638V1886:std_logic_vector(8 downto 0);
signal V254C639,V308C639,V941C639,V1041C639,V1791C639,V1887C639,C639V254,C639V308,C639V941,C639V1041,C639V1791,C639V1887:std_logic_vector(8 downto 0);
signal V255C640,V309C640,V942C640,V1042C640,V1792C640,V1888C640,C640V255,C640V309,C640V942,C640V1042,C640V1792,C640V1888:std_logic_vector(8 downto 0);
signal V256C641,V310C641,V943C641,V1043C641,V1793C641,V1889C641,C641V256,C641V310,C641V943,C641V1043,C641V1793,C641V1889:std_logic_vector(8 downto 0);
signal V257C642,V311C642,V944C642,V1044C642,V1794C642,V1890C642,C642V257,C642V311,C642V944,C642V1044,C642V1794,C642V1890:std_logic_vector(8 downto 0);
signal V258C643,V312C643,V945C643,V1045C643,V1795C643,V1891C643,C643V258,C643V312,C643V945,C643V1045,C643V1795,C643V1891:std_logic_vector(8 downto 0);
signal V259C644,V313C644,V946C644,V1046C644,V1796C644,V1892C644,C644V259,C644V313,C644V946,C644V1046,C644V1796,C644V1892:std_logic_vector(8 downto 0);
signal V260C645,V314C645,V947C645,V1047C645,V1797C645,V1893C645,C645V260,C645V314,C645V947,C645V1047,C645V1797,C645V1893:std_logic_vector(8 downto 0);
signal V261C646,V315C646,V948C646,V1048C646,V1798C646,V1894C646,C646V261,C646V315,C646V948,C646V1048,C646V1798,C646V1894:std_logic_vector(8 downto 0);
signal V262C647,V316C647,V949C647,V1049C647,V1799C647,V1895C647,C647V262,C647V316,C647V949,C647V1049,C647V1799,C647V1895:std_logic_vector(8 downto 0);
signal V263C648,V317C648,V950C648,V1050C648,V1800C648,V1896C648,C648V263,C648V317,C648V950,C648V1050,C648V1800,C648V1896:std_logic_vector(8 downto 0);
signal V264C649,V318C649,V951C649,V1051C649,V1801C649,V1897C649,C649V264,C649V318,C649V951,C649V1051,C649V1801,C649V1897:std_logic_vector(8 downto 0);
signal V265C650,V319C650,V952C650,V1052C650,V1802C650,V1898C650,C650V265,C650V319,C650V952,C650V1052,C650V1802,C650V1898:std_logic_vector(8 downto 0);
signal V266C651,V320C651,V953C651,V1053C651,V1803C651,V1899C651,C651V266,C651V320,C651V953,C651V1053,C651V1803,C651V1899:std_logic_vector(8 downto 0);
signal V267C652,V321C652,V954C652,V1054C652,V1804C652,V1900C652,C652V267,C652V321,C652V954,C652V1054,C652V1804,C652V1900:std_logic_vector(8 downto 0);
signal V268C653,V322C653,V955C653,V1055C653,V1805C653,V1901C653,C653V268,C653V322,C653V955,C653V1055,C653V1805,C653V1901:std_logic_vector(8 downto 0);
signal V269C654,V323C654,V956C654,V1056C654,V1806C654,V1902C654,C654V269,C654V323,C654V956,C654V1056,C654V1806,C654V1902:std_logic_vector(8 downto 0);
signal V270C655,V324C655,V957C655,V961C655,V1807C655,V1903C655,C655V270,C655V324,C655V957,C655V961,C655V1807,C655V1903:std_logic_vector(8 downto 0);
signal V271C656,V325C656,V958C656,V962C656,V1808C656,V1904C656,C656V271,C656V325,C656V958,C656V962,C656V1808,C656V1904:std_logic_vector(8 downto 0);
signal V272C657,V326C657,V959C657,V963C657,V1809C657,V1905C657,C657V272,C657V326,C657V959,C657V963,C657V1809,C657V1905:std_logic_vector(8 downto 0);
signal V273C658,V327C658,V960C658,V964C658,V1810C658,V1906C658,C658V273,C658V327,C658V960,C658V964,C658V1810,C658V1906:std_logic_vector(8 downto 0);
signal V274C659,V328C659,V865C659,V965C659,V1811C659,V1907C659,C659V274,C659V328,C659V865,C659V965,C659V1811,C659V1907:std_logic_vector(8 downto 0);
signal V275C660,V329C660,V866C660,V966C660,V1812C660,V1908C660,C660V275,C660V329,C660V866,C660V966,C660V1812,C660V1908:std_logic_vector(8 downto 0);
signal V276C661,V330C661,V867C661,V967C661,V1813C661,V1909C661,C661V276,C661V330,C661V867,C661V967,C661V1813,C661V1909:std_logic_vector(8 downto 0);
signal V277C662,V331C662,V868C662,V968C662,V1814C662,V1910C662,C662V277,C662V331,C662V868,C662V968,C662V1814,C662V1910:std_logic_vector(8 downto 0);
signal V278C663,V332C663,V869C663,V969C663,V1815C663,V1911C663,C663V278,C663V332,C663V869,C663V969,C663V1815,C663V1911:std_logic_vector(8 downto 0);
signal V279C664,V333C664,V870C664,V970C664,V1816C664,V1912C664,C664V279,C664V333,C664V870,C664V970,C664V1816,C664V1912:std_logic_vector(8 downto 0);
signal V280C665,V334C665,V871C665,V971C665,V1817C665,V1913C665,C665V280,C665V334,C665V871,C665V971,C665V1817,C665V1913:std_logic_vector(8 downto 0);
signal V281C666,V335C666,V872C666,V972C666,V1818C666,V1914C666,C666V281,C666V335,C666V872,C666V972,C666V1818,C666V1914:std_logic_vector(8 downto 0);
signal V282C667,V336C667,V873C667,V973C667,V1819C667,V1915C667,C667V282,C667V336,C667V873,C667V973,C667V1819,C667V1915:std_logic_vector(8 downto 0);
signal V283C668,V337C668,V874C668,V974C668,V1820C668,V1916C668,C668V283,C668V337,C668V874,C668V974,C668V1820,C668V1916:std_logic_vector(8 downto 0);
signal V284C669,V338C669,V875C669,V975C669,V1821C669,V1917C669,C669V284,C669V338,C669V875,C669V975,C669V1821,C669V1917:std_logic_vector(8 downto 0);
signal V285C670,V339C670,V876C670,V976C670,V1822C670,V1918C670,C670V285,C670V339,C670V876,C670V976,C670V1822,C670V1918:std_logic_vector(8 downto 0);
signal V286C671,V340C671,V877C671,V977C671,V1823C671,V1919C671,C671V286,C671V340,C671V877,C671V977,C671V1823,C671V1919:std_logic_vector(8 downto 0);
signal V287C672,V341C672,V878C672,V978C672,V1824C672,V1920C672,C672V287,C672V341,C672V878,C672V978,C672V1824,C672V1920:std_logic_vector(8 downto 0);
signal V108C673,V266C673,V579C673,V912C673,V1825C673,V1921C673,C673V108,C673V266,C673V579,C673V912,C673V1825,C673V1921:std_logic_vector(8 downto 0);
signal V109C674,V267C674,V580C674,V913C674,V1826C674,V1922C674,C674V109,C674V267,C674V580,C674V913,C674V1826,C674V1922:std_logic_vector(8 downto 0);
signal V110C675,V268C675,V581C675,V914C675,V1827C675,V1923C675,C675V110,C675V268,C675V581,C675V914,C675V1827,C675V1923:std_logic_vector(8 downto 0);
signal V111C676,V269C676,V582C676,V915C676,V1828C676,V1924C676,C676V111,C676V269,C676V582,C676V915,C676V1828,C676V1924:std_logic_vector(8 downto 0);
signal V112C677,V270C677,V583C677,V916C677,V1829C677,V1925C677,C677V112,C677V270,C677V583,C677V916,C677V1829,C677V1925:std_logic_vector(8 downto 0);
signal V113C678,V271C678,V584C678,V917C678,V1830C678,V1926C678,C678V113,C678V271,C678V584,C678V917,C678V1830,C678V1926:std_logic_vector(8 downto 0);
signal V114C679,V272C679,V585C679,V918C679,V1831C679,V1927C679,C679V114,C679V272,C679V585,C679V918,C679V1831,C679V1927:std_logic_vector(8 downto 0);
signal V115C680,V273C680,V586C680,V919C680,V1832C680,V1928C680,C680V115,C680V273,C680V586,C680V919,C680V1832,C680V1928:std_logic_vector(8 downto 0);
signal V116C681,V274C681,V587C681,V920C681,V1833C681,V1929C681,C681V116,C681V274,C681V587,C681V920,C681V1833,C681V1929:std_logic_vector(8 downto 0);
signal V117C682,V275C682,V588C682,V921C682,V1834C682,V1930C682,C682V117,C682V275,C682V588,C682V921,C682V1834,C682V1930:std_logic_vector(8 downto 0);
signal V118C683,V276C683,V589C683,V922C683,V1835C683,V1931C683,C683V118,C683V276,C683V589,C683V922,C683V1835,C683V1931:std_logic_vector(8 downto 0);
signal V119C684,V277C684,V590C684,V923C684,V1836C684,V1932C684,C684V119,C684V277,C684V590,C684V923,C684V1836,C684V1932:std_logic_vector(8 downto 0);
signal V120C685,V278C685,V591C685,V924C685,V1837C685,V1933C685,C685V120,C685V278,C685V591,C685V924,C685V1837,C685V1933:std_logic_vector(8 downto 0);
signal V121C686,V279C686,V592C686,V925C686,V1838C686,V1934C686,C686V121,C686V279,C686V592,C686V925,C686V1838,C686V1934:std_logic_vector(8 downto 0);
signal V122C687,V280C687,V593C687,V926C687,V1839C687,V1935C687,C687V122,C687V280,C687V593,C687V926,C687V1839,C687V1935:std_logic_vector(8 downto 0);
signal V123C688,V281C688,V594C688,V927C688,V1840C688,V1936C688,C688V123,C688V281,C688V594,C688V927,C688V1840,C688V1936:std_logic_vector(8 downto 0);
signal V124C689,V282C689,V595C689,V928C689,V1841C689,V1937C689,C689V124,C689V282,C689V595,C689V928,C689V1841,C689V1937:std_logic_vector(8 downto 0);
signal V125C690,V283C690,V596C690,V929C690,V1842C690,V1938C690,C690V125,C690V283,C690V596,C690V929,C690V1842,C690V1938:std_logic_vector(8 downto 0);
signal V126C691,V284C691,V597C691,V930C691,V1843C691,V1939C691,C691V126,C691V284,C691V597,C691V930,C691V1843,C691V1939:std_logic_vector(8 downto 0);
signal V127C692,V285C692,V598C692,V931C692,V1844C692,V1940C692,C692V127,C692V285,C692V598,C692V931,C692V1844,C692V1940:std_logic_vector(8 downto 0);
signal V128C693,V286C693,V599C693,V932C693,V1845C693,V1941C693,C693V128,C693V286,C693V599,C693V932,C693V1845,C693V1941:std_logic_vector(8 downto 0);
signal V129C694,V287C694,V600C694,V933C694,V1846C694,V1942C694,C694V129,C694V287,C694V600,C694V933,C694V1846,C694V1942:std_logic_vector(8 downto 0);
signal V130C695,V288C695,V601C695,V934C695,V1847C695,V1943C695,C695V130,C695V288,C695V601,C695V934,C695V1847,C695V1943:std_logic_vector(8 downto 0);
signal V131C696,V193C696,V602C696,V935C696,V1848C696,V1944C696,C696V131,C696V193,C696V602,C696V935,C696V1848,C696V1944:std_logic_vector(8 downto 0);
signal V132C697,V194C697,V603C697,V936C697,V1849C697,V1945C697,C697V132,C697V194,C697V603,C697V936,C697V1849,C697V1945:std_logic_vector(8 downto 0);
signal V133C698,V195C698,V604C698,V937C698,V1850C698,V1946C698,C698V133,C698V195,C698V604,C698V937,C698V1850,C698V1946:std_logic_vector(8 downto 0);
signal V134C699,V196C699,V605C699,V938C699,V1851C699,V1947C699,C699V134,C699V196,C699V605,C699V938,C699V1851,C699V1947:std_logic_vector(8 downto 0);
signal V135C700,V197C700,V606C700,V939C700,V1852C700,V1948C700,C700V135,C700V197,C700V606,C700V939,C700V1852,C700V1948:std_logic_vector(8 downto 0);
signal V136C701,V198C701,V607C701,V940C701,V1853C701,V1949C701,C701V136,C701V198,C701V607,C701V940,C701V1853,C701V1949:std_logic_vector(8 downto 0);
signal V137C702,V199C702,V608C702,V941C702,V1854C702,V1950C702,C702V137,C702V199,C702V608,C702V941,C702V1854,C702V1950:std_logic_vector(8 downto 0);
signal V138C703,V200C703,V609C703,V942C703,V1855C703,V1951C703,C703V138,C703V200,C703V609,C703V942,C703V1855,C703V1951:std_logic_vector(8 downto 0);
signal V139C704,V201C704,V610C704,V943C704,V1856C704,V1952C704,C704V139,C704V201,C704V610,C704V943,C704V1856,C704V1952:std_logic_vector(8 downto 0);
signal V140C705,V202C705,V611C705,V944C705,V1857C705,V1953C705,C705V140,C705V202,C705V611,C705V944,C705V1857,C705V1953:std_logic_vector(8 downto 0);
signal V141C706,V203C706,V612C706,V945C706,V1858C706,V1954C706,C706V141,C706V203,C706V612,C706V945,C706V1858,C706V1954:std_logic_vector(8 downto 0);
signal V142C707,V204C707,V613C707,V946C707,V1859C707,V1955C707,C707V142,C707V204,C707V613,C707V946,C707V1859,C707V1955:std_logic_vector(8 downto 0);
signal V143C708,V205C708,V614C708,V947C708,V1860C708,V1956C708,C708V143,C708V205,C708V614,C708V947,C708V1860,C708V1956:std_logic_vector(8 downto 0);
signal V144C709,V206C709,V615C709,V948C709,V1861C709,V1957C709,C709V144,C709V206,C709V615,C709V948,C709V1861,C709V1957:std_logic_vector(8 downto 0);
signal V145C710,V207C710,V616C710,V949C710,V1862C710,V1958C710,C710V145,C710V207,C710V616,C710V949,C710V1862,C710V1958:std_logic_vector(8 downto 0);
signal V146C711,V208C711,V617C711,V950C711,V1863C711,V1959C711,C711V146,C711V208,C711V617,C711V950,C711V1863,C711V1959:std_logic_vector(8 downto 0);
signal V147C712,V209C712,V618C712,V951C712,V1864C712,V1960C712,C712V147,C712V209,C712V618,C712V951,C712V1864,C712V1960:std_logic_vector(8 downto 0);
signal V148C713,V210C713,V619C713,V952C713,V1865C713,V1961C713,C713V148,C713V210,C713V619,C713V952,C713V1865,C713V1961:std_logic_vector(8 downto 0);
signal V149C714,V211C714,V620C714,V953C714,V1866C714,V1962C714,C714V149,C714V211,C714V620,C714V953,C714V1866,C714V1962:std_logic_vector(8 downto 0);
signal V150C715,V212C715,V621C715,V954C715,V1867C715,V1963C715,C715V150,C715V212,C715V621,C715V954,C715V1867,C715V1963:std_logic_vector(8 downto 0);
signal V151C716,V213C716,V622C716,V955C716,V1868C716,V1964C716,C716V151,C716V213,C716V622,C716V955,C716V1868,C716V1964:std_logic_vector(8 downto 0);
signal V152C717,V214C717,V623C717,V956C717,V1869C717,V1965C717,C717V152,C717V214,C717V623,C717V956,C717V1869,C717V1965:std_logic_vector(8 downto 0);
signal V153C718,V215C718,V624C718,V957C718,V1870C718,V1966C718,C718V153,C718V215,C718V624,C718V957,C718V1870,C718V1966:std_logic_vector(8 downto 0);
signal V154C719,V216C719,V625C719,V958C719,V1871C719,V1967C719,C719V154,C719V216,C719V625,C719V958,C719V1871,C719V1967:std_logic_vector(8 downto 0);
signal V155C720,V217C720,V626C720,V959C720,V1872C720,V1968C720,C720V155,C720V217,C720V626,C720V959,C720V1872,C720V1968:std_logic_vector(8 downto 0);
signal V156C721,V218C721,V627C721,V960C721,V1873C721,V1969C721,C721V156,C721V218,C721V627,C721V960,C721V1873,C721V1969:std_logic_vector(8 downto 0);
signal V157C722,V219C722,V628C722,V865C722,V1874C722,V1970C722,C722V157,C722V219,C722V628,C722V865,C722V1874,C722V1970:std_logic_vector(8 downto 0);
signal V158C723,V220C723,V629C723,V866C723,V1875C723,V1971C723,C723V158,C723V220,C723V629,C723V866,C723V1875,C723V1971:std_logic_vector(8 downto 0);
signal V159C724,V221C724,V630C724,V867C724,V1876C724,V1972C724,C724V159,C724V221,C724V630,C724V867,C724V1876,C724V1972:std_logic_vector(8 downto 0);
signal V160C725,V222C725,V631C725,V868C725,V1877C725,V1973C725,C725V160,C725V222,C725V631,C725V868,C725V1877,C725V1973:std_logic_vector(8 downto 0);
signal V161C726,V223C726,V632C726,V869C726,V1878C726,V1974C726,C726V161,C726V223,C726V632,C726V869,C726V1878,C726V1974:std_logic_vector(8 downto 0);
signal V162C727,V224C727,V633C727,V870C727,V1879C727,V1975C727,C727V162,C727V224,C727V633,C727V870,C727V1879,C727V1975:std_logic_vector(8 downto 0);
signal V163C728,V225C728,V634C728,V871C728,V1880C728,V1976C728,C728V163,C728V225,C728V634,C728V871,C728V1880,C728V1976:std_logic_vector(8 downto 0);
signal V164C729,V226C729,V635C729,V872C729,V1881C729,V1977C729,C729V164,C729V226,C729V635,C729V872,C729V1881,C729V1977:std_logic_vector(8 downto 0);
signal V165C730,V227C730,V636C730,V873C730,V1882C730,V1978C730,C730V165,C730V227,C730V636,C730V873,C730V1882,C730V1978:std_logic_vector(8 downto 0);
signal V166C731,V228C731,V637C731,V874C731,V1883C731,V1979C731,C731V166,C731V228,C731V637,C731V874,C731V1883,C731V1979:std_logic_vector(8 downto 0);
signal V167C732,V229C732,V638C732,V875C732,V1884C732,V1980C732,C732V167,C732V229,C732V638,C732V875,C732V1884,C732V1980:std_logic_vector(8 downto 0);
signal V168C733,V230C733,V639C733,V876C733,V1885C733,V1981C733,C733V168,C733V230,C733V639,C733V876,C733V1885,C733V1981:std_logic_vector(8 downto 0);
signal V169C734,V231C734,V640C734,V877C734,V1886C734,V1982C734,C734V169,C734V231,C734V640,C734V877,C734V1886,C734V1982:std_logic_vector(8 downto 0);
signal V170C735,V232C735,V641C735,V878C735,V1887C735,V1983C735,C735V170,C735V232,C735V641,C735V878,C735V1887,C735V1983:std_logic_vector(8 downto 0);
signal V171C736,V233C736,V642C736,V879C736,V1888C736,V1984C736,C736V171,C736V233,C736V642,C736V879,C736V1888,C736V1984:std_logic_vector(8 downto 0);
signal V172C737,V234C737,V643C737,V880C737,V1889C737,V1985C737,C737V172,C737V234,C737V643,C737V880,C737V1889,C737V1985:std_logic_vector(8 downto 0);
signal V173C738,V235C738,V644C738,V881C738,V1890C738,V1986C738,C738V173,C738V235,C738V644,C738V881,C738V1890,C738V1986:std_logic_vector(8 downto 0);
signal V174C739,V236C739,V645C739,V882C739,V1891C739,V1987C739,C739V174,C739V236,C739V645,C739V882,C739V1891,C739V1987:std_logic_vector(8 downto 0);
signal V175C740,V237C740,V646C740,V883C740,V1892C740,V1988C740,C740V175,C740V237,C740V646,C740V883,C740V1892,C740V1988:std_logic_vector(8 downto 0);
signal V176C741,V238C741,V647C741,V884C741,V1893C741,V1989C741,C741V176,C741V238,C741V647,C741V884,C741V1893,C741V1989:std_logic_vector(8 downto 0);
signal V177C742,V239C742,V648C742,V885C742,V1894C742,V1990C742,C742V177,C742V239,C742V648,C742V885,C742V1894,C742V1990:std_logic_vector(8 downto 0);
signal V178C743,V240C743,V649C743,V886C743,V1895C743,V1991C743,C743V178,C743V240,C743V649,C743V886,C743V1895,C743V1991:std_logic_vector(8 downto 0);
signal V179C744,V241C744,V650C744,V887C744,V1896C744,V1992C744,C744V179,C744V241,C744V650,C744V887,C744V1896,C744V1992:std_logic_vector(8 downto 0);
signal V180C745,V242C745,V651C745,V888C745,V1897C745,V1993C745,C745V180,C745V242,C745V651,C745V888,C745V1897,C745V1993:std_logic_vector(8 downto 0);
signal V181C746,V243C746,V652C746,V889C746,V1898C746,V1994C746,C746V181,C746V243,C746V652,C746V889,C746V1898,C746V1994:std_logic_vector(8 downto 0);
signal V182C747,V244C747,V653C747,V890C747,V1899C747,V1995C747,C747V182,C747V244,C747V653,C747V890,C747V1899,C747V1995:std_logic_vector(8 downto 0);
signal V183C748,V245C748,V654C748,V891C748,V1900C748,V1996C748,C748V183,C748V245,C748V654,C748V891,C748V1900,C748V1996:std_logic_vector(8 downto 0);
signal V184C749,V246C749,V655C749,V892C749,V1901C749,V1997C749,C749V184,C749V246,C749V655,C749V892,C749V1901,C749V1997:std_logic_vector(8 downto 0);
signal V185C750,V247C750,V656C750,V893C750,V1902C750,V1998C750,C750V185,C750V247,C750V656,C750V893,C750V1902,C750V1998:std_logic_vector(8 downto 0);
signal V186C751,V248C751,V657C751,V894C751,V1903C751,V1999C751,C751V186,C751V248,C751V657,C751V894,C751V1903,C751V1999:std_logic_vector(8 downto 0);
signal V187C752,V249C752,V658C752,V895C752,V1904C752,V2000C752,C752V187,C752V249,C752V658,C752V895,C752V1904,C752V2000:std_logic_vector(8 downto 0);
signal V188C753,V250C753,V659C753,V896C753,V1905C753,V2001C753,C753V188,C753V250,C753V659,C753V896,C753V1905,C753V2001:std_logic_vector(8 downto 0);
signal V189C754,V251C754,V660C754,V897C754,V1906C754,V2002C754,C754V189,C754V251,C754V660,C754V897,C754V1906,C754V2002:std_logic_vector(8 downto 0);
signal V190C755,V252C755,V661C755,V898C755,V1907C755,V2003C755,C755V190,C755V252,C755V661,C755V898,C755V1907,C755V2003:std_logic_vector(8 downto 0);
signal V191C756,V253C756,V662C756,V899C756,V1908C756,V2004C756,C756V191,C756V253,C756V662,C756V899,C756V1908,C756V2004:std_logic_vector(8 downto 0);
signal V192C757,V254C757,V663C757,V900C757,V1909C757,V2005C757,C757V192,C757V254,C757V663,C757V900,C757V1909,C757V2005:std_logic_vector(8 downto 0);
signal V97C758,V255C758,V664C758,V901C758,V1910C758,V2006C758,C758V97,C758V255,C758V664,C758V901,C758V1910,C758V2006:std_logic_vector(8 downto 0);
signal V98C759,V256C759,V665C759,V902C759,V1911C759,V2007C759,C759V98,C759V256,C759V665,C759V902,C759V1911,C759V2007:std_logic_vector(8 downto 0);
signal V99C760,V257C760,V666C760,V903C760,V1912C760,V2008C760,C760V99,C760V257,C760V666,C760V903,C760V1912,C760V2008:std_logic_vector(8 downto 0);
signal V100C761,V258C761,V667C761,V904C761,V1913C761,V2009C761,C761V100,C761V258,C761V667,C761V904,C761V1913,C761V2009:std_logic_vector(8 downto 0);
signal V101C762,V259C762,V668C762,V905C762,V1914C762,V2010C762,C762V101,C762V259,C762V668,C762V905,C762V1914,C762V2010:std_logic_vector(8 downto 0);
signal V102C763,V260C763,V669C763,V906C763,V1915C763,V2011C763,C763V102,C763V260,C763V669,C763V906,C763V1915,C763V2011:std_logic_vector(8 downto 0);
signal V103C764,V261C764,V670C764,V907C764,V1916C764,V2012C764,C764V103,C764V261,C764V670,C764V907,C764V1916,C764V2012:std_logic_vector(8 downto 0);
signal V104C765,V262C765,V671C765,V908C765,V1917C765,V2013C765,C765V104,C765V262,C765V671,C765V908,C765V1917,C765V2013:std_logic_vector(8 downto 0);
signal V105C766,V263C766,V672C766,V909C766,V1918C766,V2014C766,C766V105,C766V263,C766V672,C766V909,C766V1918,C766V2014:std_logic_vector(8 downto 0);
signal V106C767,V264C767,V577C767,V910C767,V1919C767,V2015C767,C767V106,C767V264,C767V577,C767V910,C767V1919,C767V2015:std_logic_vector(8 downto 0);
signal V107C768,V265C768,V578C768,V911C768,V1920C768,V2016C768,C768V107,C768V265,C768V578,C768V911,C768V1920,C768V2016:std_logic_vector(8 downto 0);
signal V13C769,V468C769,V505C769,V716C769,V1108C769,V1921C769,V2017C769,C769V13,C769V468,C769V505,C769V716,C769V1108,C769V1921,C769V2017:std_logic_vector(8 downto 0);
signal V14C770,V469C770,V506C770,V717C770,V1109C770,V1922C770,V2018C770,C770V14,C770V469,C770V506,C770V717,C770V1109,C770V1922,C770V2018:std_logic_vector(8 downto 0);
signal V15C771,V470C771,V507C771,V718C771,V1110C771,V1923C771,V2019C771,C771V15,C771V470,C771V507,C771V718,C771V1110,C771V1923,C771V2019:std_logic_vector(8 downto 0);
signal V16C772,V471C772,V508C772,V719C772,V1111C772,V1924C772,V2020C772,C772V16,C772V471,C772V508,C772V719,C772V1111,C772V1924,C772V2020:std_logic_vector(8 downto 0);
signal V17C773,V472C773,V509C773,V720C773,V1112C773,V1925C773,V2021C773,C773V17,C773V472,C773V509,C773V720,C773V1112,C773V1925,C773V2021:std_logic_vector(8 downto 0);
signal V18C774,V473C774,V510C774,V721C774,V1113C774,V1926C774,V2022C774,C774V18,C774V473,C774V510,C774V721,C774V1113,C774V1926,C774V2022:std_logic_vector(8 downto 0);
signal V19C775,V474C775,V511C775,V722C775,V1114C775,V1927C775,V2023C775,C775V19,C775V474,C775V511,C775V722,C775V1114,C775V1927,C775V2023:std_logic_vector(8 downto 0);
signal V20C776,V475C776,V512C776,V723C776,V1115C776,V1928C776,V2024C776,C776V20,C776V475,C776V512,C776V723,C776V1115,C776V1928,C776V2024:std_logic_vector(8 downto 0);
signal V21C777,V476C777,V513C777,V724C777,V1116C777,V1929C777,V2025C777,C777V21,C777V476,C777V513,C777V724,C777V1116,C777V1929,C777V2025:std_logic_vector(8 downto 0);
signal V22C778,V477C778,V514C778,V725C778,V1117C778,V1930C778,V2026C778,C778V22,C778V477,C778V514,C778V725,C778V1117,C778V1930,C778V2026:std_logic_vector(8 downto 0);
signal V23C779,V478C779,V515C779,V726C779,V1118C779,V1931C779,V2027C779,C779V23,C779V478,C779V515,C779V726,C779V1118,C779V1931,C779V2027:std_logic_vector(8 downto 0);
signal V24C780,V479C780,V516C780,V727C780,V1119C780,V1932C780,V2028C780,C780V24,C780V479,C780V516,C780V727,C780V1119,C780V1932,C780V2028:std_logic_vector(8 downto 0);
signal V25C781,V480C781,V517C781,V728C781,V1120C781,V1933C781,V2029C781,C781V25,C781V480,C781V517,C781V728,C781V1120,C781V1933,C781V2029:std_logic_vector(8 downto 0);
signal V26C782,V385C782,V518C782,V729C782,V1121C782,V1934C782,V2030C782,C782V26,C782V385,C782V518,C782V729,C782V1121,C782V1934,C782V2030:std_logic_vector(8 downto 0);
signal V27C783,V386C783,V519C783,V730C783,V1122C783,V1935C783,V2031C783,C783V27,C783V386,C783V519,C783V730,C783V1122,C783V1935,C783V2031:std_logic_vector(8 downto 0);
signal V28C784,V387C784,V520C784,V731C784,V1123C784,V1936C784,V2032C784,C784V28,C784V387,C784V520,C784V731,C784V1123,C784V1936,C784V2032:std_logic_vector(8 downto 0);
signal V29C785,V388C785,V521C785,V732C785,V1124C785,V1937C785,V2033C785,C785V29,C785V388,C785V521,C785V732,C785V1124,C785V1937,C785V2033:std_logic_vector(8 downto 0);
signal V30C786,V389C786,V522C786,V733C786,V1125C786,V1938C786,V2034C786,C786V30,C786V389,C786V522,C786V733,C786V1125,C786V1938,C786V2034:std_logic_vector(8 downto 0);
signal V31C787,V390C787,V523C787,V734C787,V1126C787,V1939C787,V2035C787,C787V31,C787V390,C787V523,C787V734,C787V1126,C787V1939,C787V2035:std_logic_vector(8 downto 0);
signal V32C788,V391C788,V524C788,V735C788,V1127C788,V1940C788,V2036C788,C788V32,C788V391,C788V524,C788V735,C788V1127,C788V1940,C788V2036:std_logic_vector(8 downto 0);
signal V33C789,V392C789,V525C789,V736C789,V1128C789,V1941C789,V2037C789,C789V33,C789V392,C789V525,C789V736,C789V1128,C789V1941,C789V2037:std_logic_vector(8 downto 0);
signal V34C790,V393C790,V526C790,V737C790,V1129C790,V1942C790,V2038C790,C790V34,C790V393,C790V526,C790V737,C790V1129,C790V1942,C790V2038:std_logic_vector(8 downto 0);
signal V35C791,V394C791,V527C791,V738C791,V1130C791,V1943C791,V2039C791,C791V35,C791V394,C791V527,C791V738,C791V1130,C791V1943,C791V2039:std_logic_vector(8 downto 0);
signal V36C792,V395C792,V528C792,V739C792,V1131C792,V1944C792,V2040C792,C792V36,C792V395,C792V528,C792V739,C792V1131,C792V1944,C792V2040:std_logic_vector(8 downto 0);
signal V37C793,V396C793,V529C793,V740C793,V1132C793,V1945C793,V2041C793,C793V37,C793V396,C793V529,C793V740,C793V1132,C793V1945,C793V2041:std_logic_vector(8 downto 0);
signal V38C794,V397C794,V530C794,V741C794,V1133C794,V1946C794,V2042C794,C794V38,C794V397,C794V530,C794V741,C794V1133,C794V1946,C794V2042:std_logic_vector(8 downto 0);
signal V39C795,V398C795,V531C795,V742C795,V1134C795,V1947C795,V2043C795,C795V39,C795V398,C795V531,C795V742,C795V1134,C795V1947,C795V2043:std_logic_vector(8 downto 0);
signal V40C796,V399C796,V532C796,V743C796,V1135C796,V1948C796,V2044C796,C796V40,C796V399,C796V532,C796V743,C796V1135,C796V1948,C796V2044:std_logic_vector(8 downto 0);
signal V41C797,V400C797,V533C797,V744C797,V1136C797,V1949C797,V2045C797,C797V41,C797V400,C797V533,C797V744,C797V1136,C797V1949,C797V2045:std_logic_vector(8 downto 0);
signal V42C798,V401C798,V534C798,V745C798,V1137C798,V1950C798,V2046C798,C798V42,C798V401,C798V534,C798V745,C798V1137,C798V1950,C798V2046:std_logic_vector(8 downto 0);
signal V43C799,V402C799,V535C799,V746C799,V1138C799,V1951C799,V2047C799,C799V43,C799V402,C799V535,C799V746,C799V1138,C799V1951,C799V2047:std_logic_vector(8 downto 0);
signal V44C800,V403C800,V536C800,V747C800,V1139C800,V1952C800,V2048C800,C800V44,C800V403,C800V536,C800V747,C800V1139,C800V1952,C800V2048:std_logic_vector(8 downto 0);
signal V45C801,V404C801,V537C801,V748C801,V1140C801,V1953C801,V2049C801,C801V45,C801V404,C801V537,C801V748,C801V1140,C801V1953,C801V2049:std_logic_vector(8 downto 0);
signal V46C802,V405C802,V538C802,V749C802,V1141C802,V1954C802,V2050C802,C802V46,C802V405,C802V538,C802V749,C802V1141,C802V1954,C802V2050:std_logic_vector(8 downto 0);
signal V47C803,V406C803,V539C803,V750C803,V1142C803,V1955C803,V2051C803,C803V47,C803V406,C803V539,C803V750,C803V1142,C803V1955,C803V2051:std_logic_vector(8 downto 0);
signal V48C804,V407C804,V540C804,V751C804,V1143C804,V1956C804,V2052C804,C804V48,C804V407,C804V540,C804V751,C804V1143,C804V1956,C804V2052:std_logic_vector(8 downto 0);
signal V49C805,V408C805,V541C805,V752C805,V1144C805,V1957C805,V2053C805,C805V49,C805V408,C805V541,C805V752,C805V1144,C805V1957,C805V2053:std_logic_vector(8 downto 0);
signal V50C806,V409C806,V542C806,V753C806,V1145C806,V1958C806,V2054C806,C806V50,C806V409,C806V542,C806V753,C806V1145,C806V1958,C806V2054:std_logic_vector(8 downto 0);
signal V51C807,V410C807,V543C807,V754C807,V1146C807,V1959C807,V2055C807,C807V51,C807V410,C807V543,C807V754,C807V1146,C807V1959,C807V2055:std_logic_vector(8 downto 0);
signal V52C808,V411C808,V544C808,V755C808,V1147C808,V1960C808,V2056C808,C808V52,C808V411,C808V544,C808V755,C808V1147,C808V1960,C808V2056:std_logic_vector(8 downto 0);
signal V53C809,V412C809,V545C809,V756C809,V1148C809,V1961C809,V2057C809,C809V53,C809V412,C809V545,C809V756,C809V1148,C809V1961,C809V2057:std_logic_vector(8 downto 0);
signal V54C810,V413C810,V546C810,V757C810,V1149C810,V1962C810,V2058C810,C810V54,C810V413,C810V546,C810V757,C810V1149,C810V1962,C810V2058:std_logic_vector(8 downto 0);
signal V55C811,V414C811,V547C811,V758C811,V1150C811,V1963C811,V2059C811,C811V55,C811V414,C811V547,C811V758,C811V1150,C811V1963,C811V2059:std_logic_vector(8 downto 0);
signal V56C812,V415C812,V548C812,V759C812,V1151C812,V1964C812,V2060C812,C812V56,C812V415,C812V548,C812V759,C812V1151,C812V1964,C812V2060:std_logic_vector(8 downto 0);
signal V57C813,V416C813,V549C813,V760C813,V1152C813,V1965C813,V2061C813,C813V57,C813V416,C813V549,C813V760,C813V1152,C813V1965,C813V2061:std_logic_vector(8 downto 0);
signal V58C814,V417C814,V550C814,V761C814,V1057C814,V1966C814,V2062C814,C814V58,C814V417,C814V550,C814V761,C814V1057,C814V1966,C814V2062:std_logic_vector(8 downto 0);
signal V59C815,V418C815,V551C815,V762C815,V1058C815,V1967C815,V2063C815,C815V59,C815V418,C815V551,C815V762,C815V1058,C815V1967,C815V2063:std_logic_vector(8 downto 0);
signal V60C816,V419C816,V552C816,V763C816,V1059C816,V1968C816,V2064C816,C816V60,C816V419,C816V552,C816V763,C816V1059,C816V1968,C816V2064:std_logic_vector(8 downto 0);
signal V61C817,V420C817,V553C817,V764C817,V1060C817,V1969C817,V2065C817,C817V61,C817V420,C817V553,C817V764,C817V1060,C817V1969,C817V2065:std_logic_vector(8 downto 0);
signal V62C818,V421C818,V554C818,V765C818,V1061C818,V1970C818,V2066C818,C818V62,C818V421,C818V554,C818V765,C818V1061,C818V1970,C818V2066:std_logic_vector(8 downto 0);
signal V63C819,V422C819,V555C819,V766C819,V1062C819,V1971C819,V2067C819,C819V63,C819V422,C819V555,C819V766,C819V1062,C819V1971,C819V2067:std_logic_vector(8 downto 0);
signal V64C820,V423C820,V556C820,V767C820,V1063C820,V1972C820,V2068C820,C820V64,C820V423,C820V556,C820V767,C820V1063,C820V1972,C820V2068:std_logic_vector(8 downto 0);
signal V65C821,V424C821,V557C821,V768C821,V1064C821,V1973C821,V2069C821,C821V65,C821V424,C821V557,C821V768,C821V1064,C821V1973,C821V2069:std_logic_vector(8 downto 0);
signal V66C822,V425C822,V558C822,V673C822,V1065C822,V1974C822,V2070C822,C822V66,C822V425,C822V558,C822V673,C822V1065,C822V1974,C822V2070:std_logic_vector(8 downto 0);
signal V67C823,V426C823,V559C823,V674C823,V1066C823,V1975C823,V2071C823,C823V67,C823V426,C823V559,C823V674,C823V1066,C823V1975,C823V2071:std_logic_vector(8 downto 0);
signal V68C824,V427C824,V560C824,V675C824,V1067C824,V1976C824,V2072C824,C824V68,C824V427,C824V560,C824V675,C824V1067,C824V1976,C824V2072:std_logic_vector(8 downto 0);
signal V69C825,V428C825,V561C825,V676C825,V1068C825,V1977C825,V2073C825,C825V69,C825V428,C825V561,C825V676,C825V1068,C825V1977,C825V2073:std_logic_vector(8 downto 0);
signal V70C826,V429C826,V562C826,V677C826,V1069C826,V1978C826,V2074C826,C826V70,C826V429,C826V562,C826V677,C826V1069,C826V1978,C826V2074:std_logic_vector(8 downto 0);
signal V71C827,V430C827,V563C827,V678C827,V1070C827,V1979C827,V2075C827,C827V71,C827V430,C827V563,C827V678,C827V1070,C827V1979,C827V2075:std_logic_vector(8 downto 0);
signal V72C828,V431C828,V564C828,V679C828,V1071C828,V1980C828,V2076C828,C828V72,C828V431,C828V564,C828V679,C828V1071,C828V1980,C828V2076:std_logic_vector(8 downto 0);
signal V73C829,V432C829,V565C829,V680C829,V1072C829,V1981C829,V2077C829,C829V73,C829V432,C829V565,C829V680,C829V1072,C829V1981,C829V2077:std_logic_vector(8 downto 0);
signal V74C830,V433C830,V566C830,V681C830,V1073C830,V1982C830,V2078C830,C830V74,C830V433,C830V566,C830V681,C830V1073,C830V1982,C830V2078:std_logic_vector(8 downto 0);
signal V75C831,V434C831,V567C831,V682C831,V1074C831,V1983C831,V2079C831,C831V75,C831V434,C831V567,C831V682,C831V1074,C831V1983,C831V2079:std_logic_vector(8 downto 0);
signal V76C832,V435C832,V568C832,V683C832,V1075C832,V1984C832,V2080C832,C832V76,C832V435,C832V568,C832V683,C832V1075,C832V1984,C832V2080:std_logic_vector(8 downto 0);
signal V77C833,V436C833,V569C833,V684C833,V1076C833,V1985C833,V2081C833,C833V77,C833V436,C833V569,C833V684,C833V1076,C833V1985,C833V2081:std_logic_vector(8 downto 0);
signal V78C834,V437C834,V570C834,V685C834,V1077C834,V1986C834,V2082C834,C834V78,C834V437,C834V570,C834V685,C834V1077,C834V1986,C834V2082:std_logic_vector(8 downto 0);
signal V79C835,V438C835,V571C835,V686C835,V1078C835,V1987C835,V2083C835,C835V79,C835V438,C835V571,C835V686,C835V1078,C835V1987,C835V2083:std_logic_vector(8 downto 0);
signal V80C836,V439C836,V572C836,V687C836,V1079C836,V1988C836,V2084C836,C836V80,C836V439,C836V572,C836V687,C836V1079,C836V1988,C836V2084:std_logic_vector(8 downto 0);
signal V81C837,V440C837,V573C837,V688C837,V1080C837,V1989C837,V2085C837,C837V81,C837V440,C837V573,C837V688,C837V1080,C837V1989,C837V2085:std_logic_vector(8 downto 0);
signal V82C838,V441C838,V574C838,V689C838,V1081C838,V1990C838,V2086C838,C838V82,C838V441,C838V574,C838V689,C838V1081,C838V1990,C838V2086:std_logic_vector(8 downto 0);
signal V83C839,V442C839,V575C839,V690C839,V1082C839,V1991C839,V2087C839,C839V83,C839V442,C839V575,C839V690,C839V1082,C839V1991,C839V2087:std_logic_vector(8 downto 0);
signal V84C840,V443C840,V576C840,V691C840,V1083C840,V1992C840,V2088C840,C840V84,C840V443,C840V576,C840V691,C840V1083,C840V1992,C840V2088:std_logic_vector(8 downto 0);
signal V85C841,V444C841,V481C841,V692C841,V1084C841,V1993C841,V2089C841,C841V85,C841V444,C841V481,C841V692,C841V1084,C841V1993,C841V2089:std_logic_vector(8 downto 0);
signal V86C842,V445C842,V482C842,V693C842,V1085C842,V1994C842,V2090C842,C842V86,C842V445,C842V482,C842V693,C842V1085,C842V1994,C842V2090:std_logic_vector(8 downto 0);
signal V87C843,V446C843,V483C843,V694C843,V1086C843,V1995C843,V2091C843,C843V87,C843V446,C843V483,C843V694,C843V1086,C843V1995,C843V2091:std_logic_vector(8 downto 0);
signal V88C844,V447C844,V484C844,V695C844,V1087C844,V1996C844,V2092C844,C844V88,C844V447,C844V484,C844V695,C844V1087,C844V1996,C844V2092:std_logic_vector(8 downto 0);
signal V89C845,V448C845,V485C845,V696C845,V1088C845,V1997C845,V2093C845,C845V89,C845V448,C845V485,C845V696,C845V1088,C845V1997,C845V2093:std_logic_vector(8 downto 0);
signal V90C846,V449C846,V486C846,V697C846,V1089C846,V1998C846,V2094C846,C846V90,C846V449,C846V486,C846V697,C846V1089,C846V1998,C846V2094:std_logic_vector(8 downto 0);
signal V91C847,V450C847,V487C847,V698C847,V1090C847,V1999C847,V2095C847,C847V91,C847V450,C847V487,C847V698,C847V1090,C847V1999,C847V2095:std_logic_vector(8 downto 0);
signal V92C848,V451C848,V488C848,V699C848,V1091C848,V2000C848,V2096C848,C848V92,C848V451,C848V488,C848V699,C848V1091,C848V2000,C848V2096:std_logic_vector(8 downto 0);
signal V93C849,V452C849,V489C849,V700C849,V1092C849,V2001C849,V2097C849,C849V93,C849V452,C849V489,C849V700,C849V1092,C849V2001,C849V2097:std_logic_vector(8 downto 0);
signal V94C850,V453C850,V490C850,V701C850,V1093C850,V2002C850,V2098C850,C850V94,C850V453,C850V490,C850V701,C850V1093,C850V2002,C850V2098:std_logic_vector(8 downto 0);
signal V95C851,V454C851,V491C851,V702C851,V1094C851,V2003C851,V2099C851,C851V95,C851V454,C851V491,C851V702,C851V1094,C851V2003,C851V2099:std_logic_vector(8 downto 0);
signal V96C852,V455C852,V492C852,V703C852,V1095C852,V2004C852,V2100C852,C852V96,C852V455,C852V492,C852V703,C852V1095,C852V2004,C852V2100:std_logic_vector(8 downto 0);
signal V1C853,V456C853,V493C853,V704C853,V1096C853,V2005C853,V2101C853,C853V1,C853V456,C853V493,C853V704,C853V1096,C853V2005,C853V2101:std_logic_vector(8 downto 0);
signal V2C854,V457C854,V494C854,V705C854,V1097C854,V2006C854,V2102C854,C854V2,C854V457,C854V494,C854V705,C854V1097,C854V2006,C854V2102:std_logic_vector(8 downto 0);
signal V3C855,V458C855,V495C855,V706C855,V1098C855,V2007C855,V2103C855,C855V3,C855V458,C855V495,C855V706,C855V1098,C855V2007,C855V2103:std_logic_vector(8 downto 0);
signal V4C856,V459C856,V496C856,V707C856,V1099C856,V2008C856,V2104C856,C856V4,C856V459,C856V496,C856V707,C856V1099,C856V2008,C856V2104:std_logic_vector(8 downto 0);
signal V5C857,V460C857,V497C857,V708C857,V1100C857,V2009C857,V2105C857,C857V5,C857V460,C857V497,C857V708,C857V1100,C857V2009,C857V2105:std_logic_vector(8 downto 0);
signal V6C858,V461C858,V498C858,V709C858,V1101C858,V2010C858,V2106C858,C858V6,C858V461,C858V498,C858V709,C858V1101,C858V2010,C858V2106:std_logic_vector(8 downto 0);
signal V7C859,V462C859,V499C859,V710C859,V1102C859,V2011C859,V2107C859,C859V7,C859V462,C859V499,C859V710,C859V1102,C859V2011,C859V2107:std_logic_vector(8 downto 0);
signal V8C860,V463C860,V500C860,V711C860,V1103C860,V2012C860,V2108C860,C860V8,C860V463,C860V500,C860V711,C860V1103,C860V2012,C860V2108:std_logic_vector(8 downto 0);
signal V9C861,V464C861,V501C861,V712C861,V1104C861,V2013C861,V2109C861,C861V9,C861V464,C861V501,C861V712,C861V1104,C861V2013,C861V2109:std_logic_vector(8 downto 0);
signal V10C862,V465C862,V502C862,V713C862,V1105C862,V2014C862,V2110C862,C862V10,C862V465,C862V502,C862V713,C862V1105,C862V2014,C862V2110:std_logic_vector(8 downto 0);
signal V11C863,V466C863,V503C863,V714C863,V1106C863,V2015C863,V2111C863,C863V11,C863V466,C863V503,C863V714,C863V1106,C863V2015,C863V2111:std_logic_vector(8 downto 0);
signal V12C864,V467C864,V504C864,V715C864,V1107C864,V2016C864,V2112C864,C864V12,C864V467,C864V504,C864V715,C864V1107,C864V2016,C864V2112:std_logic_vector(8 downto 0);
signal V575C865,V732C865,V1031C865,V1129C865,V2017C865,V2113C865,C865V575,C865V732,C865V1031,C865V1129,C865V2017,C865V2113:std_logic_vector(8 downto 0);
signal V576C866,V733C866,V1032C866,V1130C866,V2018C866,V2114C866,C866V576,C866V733,C866V1032,C866V1130,C866V2018,C866V2114:std_logic_vector(8 downto 0);
signal V481C867,V734C867,V1033C867,V1131C867,V2019C867,V2115C867,C867V481,C867V734,C867V1033,C867V1131,C867V2019,C867V2115:std_logic_vector(8 downto 0);
signal V482C868,V735C868,V1034C868,V1132C868,V2020C868,V2116C868,C868V482,C868V735,C868V1034,C868V1132,C868V2020,C868V2116:std_logic_vector(8 downto 0);
signal V483C869,V736C869,V1035C869,V1133C869,V2021C869,V2117C869,C869V483,C869V736,C869V1035,C869V1133,C869V2021,C869V2117:std_logic_vector(8 downto 0);
signal V484C870,V737C870,V1036C870,V1134C870,V2022C870,V2118C870,C870V484,C870V737,C870V1036,C870V1134,C870V2022,C870V2118:std_logic_vector(8 downto 0);
signal V485C871,V738C871,V1037C871,V1135C871,V2023C871,V2119C871,C871V485,C871V738,C871V1037,C871V1135,C871V2023,C871V2119:std_logic_vector(8 downto 0);
signal V486C872,V739C872,V1038C872,V1136C872,V2024C872,V2120C872,C872V486,C872V739,C872V1038,C872V1136,C872V2024,C872V2120:std_logic_vector(8 downto 0);
signal V487C873,V740C873,V1039C873,V1137C873,V2025C873,V2121C873,C873V487,C873V740,C873V1039,C873V1137,C873V2025,C873V2121:std_logic_vector(8 downto 0);
signal V488C874,V741C874,V1040C874,V1138C874,V2026C874,V2122C874,C874V488,C874V741,C874V1040,C874V1138,C874V2026,C874V2122:std_logic_vector(8 downto 0);
signal V489C875,V742C875,V1041C875,V1139C875,V2027C875,V2123C875,C875V489,C875V742,C875V1041,C875V1139,C875V2027,C875V2123:std_logic_vector(8 downto 0);
signal V490C876,V743C876,V1042C876,V1140C876,V2028C876,V2124C876,C876V490,C876V743,C876V1042,C876V1140,C876V2028,C876V2124:std_logic_vector(8 downto 0);
signal V491C877,V744C877,V1043C877,V1141C877,V2029C877,V2125C877,C877V491,C877V744,C877V1043,C877V1141,C877V2029,C877V2125:std_logic_vector(8 downto 0);
signal V492C878,V745C878,V1044C878,V1142C878,V2030C878,V2126C878,C878V492,C878V745,C878V1044,C878V1142,C878V2030,C878V2126:std_logic_vector(8 downto 0);
signal V493C879,V746C879,V1045C879,V1143C879,V2031C879,V2127C879,C879V493,C879V746,C879V1045,C879V1143,C879V2031,C879V2127:std_logic_vector(8 downto 0);
signal V494C880,V747C880,V1046C880,V1144C880,V2032C880,V2128C880,C880V494,C880V747,C880V1046,C880V1144,C880V2032,C880V2128:std_logic_vector(8 downto 0);
signal V495C881,V748C881,V1047C881,V1145C881,V2033C881,V2129C881,C881V495,C881V748,C881V1047,C881V1145,C881V2033,C881V2129:std_logic_vector(8 downto 0);
signal V496C882,V749C882,V1048C882,V1146C882,V2034C882,V2130C882,C882V496,C882V749,C882V1048,C882V1146,C882V2034,C882V2130:std_logic_vector(8 downto 0);
signal V497C883,V750C883,V1049C883,V1147C883,V2035C883,V2131C883,C883V497,C883V750,C883V1049,C883V1147,C883V2035,C883V2131:std_logic_vector(8 downto 0);
signal V498C884,V751C884,V1050C884,V1148C884,V2036C884,V2132C884,C884V498,C884V751,C884V1050,C884V1148,C884V2036,C884V2132:std_logic_vector(8 downto 0);
signal V499C885,V752C885,V1051C885,V1149C885,V2037C885,V2133C885,C885V499,C885V752,C885V1051,C885V1149,C885V2037,C885V2133:std_logic_vector(8 downto 0);
signal V500C886,V753C886,V1052C886,V1150C886,V2038C886,V2134C886,C886V500,C886V753,C886V1052,C886V1150,C886V2038,C886V2134:std_logic_vector(8 downto 0);
signal V501C887,V754C887,V1053C887,V1151C887,V2039C887,V2135C887,C887V501,C887V754,C887V1053,C887V1151,C887V2039,C887V2135:std_logic_vector(8 downto 0);
signal V502C888,V755C888,V1054C888,V1152C888,V2040C888,V2136C888,C888V502,C888V755,C888V1054,C888V1152,C888V2040,C888V2136:std_logic_vector(8 downto 0);
signal V503C889,V756C889,V1055C889,V1057C889,V2041C889,V2137C889,C889V503,C889V756,C889V1055,C889V1057,C889V2041,C889V2137:std_logic_vector(8 downto 0);
signal V504C890,V757C890,V1056C890,V1058C890,V2042C890,V2138C890,C890V504,C890V757,C890V1056,C890V1058,C890V2042,C890V2138:std_logic_vector(8 downto 0);
signal V505C891,V758C891,V961C891,V1059C891,V2043C891,V2139C891,C891V505,C891V758,C891V961,C891V1059,C891V2043,C891V2139:std_logic_vector(8 downto 0);
signal V506C892,V759C892,V962C892,V1060C892,V2044C892,V2140C892,C892V506,C892V759,C892V962,C892V1060,C892V2044,C892V2140:std_logic_vector(8 downto 0);
signal V507C893,V760C893,V963C893,V1061C893,V2045C893,V2141C893,C893V507,C893V760,C893V963,C893V1061,C893V2045,C893V2141:std_logic_vector(8 downto 0);
signal V508C894,V761C894,V964C894,V1062C894,V2046C894,V2142C894,C894V508,C894V761,C894V964,C894V1062,C894V2046,C894V2142:std_logic_vector(8 downto 0);
signal V509C895,V762C895,V965C895,V1063C895,V2047C895,V2143C895,C895V509,C895V762,C895V965,C895V1063,C895V2047,C895V2143:std_logic_vector(8 downto 0);
signal V510C896,V763C896,V966C896,V1064C896,V2048C896,V2144C896,C896V510,C896V763,C896V966,C896V1064,C896V2048,C896V2144:std_logic_vector(8 downto 0);
signal V511C897,V764C897,V967C897,V1065C897,V2049C897,V2145C897,C897V511,C897V764,C897V967,C897V1065,C897V2049,C897V2145:std_logic_vector(8 downto 0);
signal V512C898,V765C898,V968C898,V1066C898,V2050C898,V2146C898,C898V512,C898V765,C898V968,C898V1066,C898V2050,C898V2146:std_logic_vector(8 downto 0);
signal V513C899,V766C899,V969C899,V1067C899,V2051C899,V2147C899,C899V513,C899V766,C899V969,C899V1067,C899V2051,C899V2147:std_logic_vector(8 downto 0);
signal V514C900,V767C900,V970C900,V1068C900,V2052C900,V2148C900,C900V514,C900V767,C900V970,C900V1068,C900V2052,C900V2148:std_logic_vector(8 downto 0);
signal V515C901,V768C901,V971C901,V1069C901,V2053C901,V2149C901,C901V515,C901V768,C901V971,C901V1069,C901V2053,C901V2149:std_logic_vector(8 downto 0);
signal V516C902,V673C902,V972C902,V1070C902,V2054C902,V2150C902,C902V516,C902V673,C902V972,C902V1070,C902V2054,C902V2150:std_logic_vector(8 downto 0);
signal V517C903,V674C903,V973C903,V1071C903,V2055C903,V2151C903,C903V517,C903V674,C903V973,C903V1071,C903V2055,C903V2151:std_logic_vector(8 downto 0);
signal V518C904,V675C904,V974C904,V1072C904,V2056C904,V2152C904,C904V518,C904V675,C904V974,C904V1072,C904V2056,C904V2152:std_logic_vector(8 downto 0);
signal V519C905,V676C905,V975C905,V1073C905,V2057C905,V2153C905,C905V519,C905V676,C905V975,C905V1073,C905V2057,C905V2153:std_logic_vector(8 downto 0);
signal V520C906,V677C906,V976C906,V1074C906,V2058C906,V2154C906,C906V520,C906V677,C906V976,C906V1074,C906V2058,C906V2154:std_logic_vector(8 downto 0);
signal V521C907,V678C907,V977C907,V1075C907,V2059C907,V2155C907,C907V521,C907V678,C907V977,C907V1075,C907V2059,C907V2155:std_logic_vector(8 downto 0);
signal V522C908,V679C908,V978C908,V1076C908,V2060C908,V2156C908,C908V522,C908V679,C908V978,C908V1076,C908V2060,C908V2156:std_logic_vector(8 downto 0);
signal V523C909,V680C909,V979C909,V1077C909,V2061C909,V2157C909,C909V523,C909V680,C909V979,C909V1077,C909V2061,C909V2157:std_logic_vector(8 downto 0);
signal V524C910,V681C910,V980C910,V1078C910,V2062C910,V2158C910,C910V524,C910V681,C910V980,C910V1078,C910V2062,C910V2158:std_logic_vector(8 downto 0);
signal V525C911,V682C911,V981C911,V1079C911,V2063C911,V2159C911,C911V525,C911V682,C911V981,C911V1079,C911V2063,C911V2159:std_logic_vector(8 downto 0);
signal V526C912,V683C912,V982C912,V1080C912,V2064C912,V2160C912,C912V526,C912V683,C912V982,C912V1080,C912V2064,C912V2160:std_logic_vector(8 downto 0);
signal V527C913,V684C913,V983C913,V1081C913,V2065C913,V2161C913,C913V527,C913V684,C913V983,C913V1081,C913V2065,C913V2161:std_logic_vector(8 downto 0);
signal V528C914,V685C914,V984C914,V1082C914,V2066C914,V2162C914,C914V528,C914V685,C914V984,C914V1082,C914V2066,C914V2162:std_logic_vector(8 downto 0);
signal V529C915,V686C915,V985C915,V1083C915,V2067C915,V2163C915,C915V529,C915V686,C915V985,C915V1083,C915V2067,C915V2163:std_logic_vector(8 downto 0);
signal V530C916,V687C916,V986C916,V1084C916,V2068C916,V2164C916,C916V530,C916V687,C916V986,C916V1084,C916V2068,C916V2164:std_logic_vector(8 downto 0);
signal V531C917,V688C917,V987C917,V1085C917,V2069C917,V2165C917,C917V531,C917V688,C917V987,C917V1085,C917V2069,C917V2165:std_logic_vector(8 downto 0);
signal V532C918,V689C918,V988C918,V1086C918,V2070C918,V2166C918,C918V532,C918V689,C918V988,C918V1086,C918V2070,C918V2166:std_logic_vector(8 downto 0);
signal V533C919,V690C919,V989C919,V1087C919,V2071C919,V2167C919,C919V533,C919V690,C919V989,C919V1087,C919V2071,C919V2167:std_logic_vector(8 downto 0);
signal V534C920,V691C920,V990C920,V1088C920,V2072C920,V2168C920,C920V534,C920V691,C920V990,C920V1088,C920V2072,C920V2168:std_logic_vector(8 downto 0);
signal V535C921,V692C921,V991C921,V1089C921,V2073C921,V2169C921,C921V535,C921V692,C921V991,C921V1089,C921V2073,C921V2169:std_logic_vector(8 downto 0);
signal V536C922,V693C922,V992C922,V1090C922,V2074C922,V2170C922,C922V536,C922V693,C922V992,C922V1090,C922V2074,C922V2170:std_logic_vector(8 downto 0);
signal V537C923,V694C923,V993C923,V1091C923,V2075C923,V2171C923,C923V537,C923V694,C923V993,C923V1091,C923V2075,C923V2171:std_logic_vector(8 downto 0);
signal V538C924,V695C924,V994C924,V1092C924,V2076C924,V2172C924,C924V538,C924V695,C924V994,C924V1092,C924V2076,C924V2172:std_logic_vector(8 downto 0);
signal V539C925,V696C925,V995C925,V1093C925,V2077C925,V2173C925,C925V539,C925V696,C925V995,C925V1093,C925V2077,C925V2173:std_logic_vector(8 downto 0);
signal V540C926,V697C926,V996C926,V1094C926,V2078C926,V2174C926,C926V540,C926V697,C926V996,C926V1094,C926V2078,C926V2174:std_logic_vector(8 downto 0);
signal V541C927,V698C927,V997C927,V1095C927,V2079C927,V2175C927,C927V541,C927V698,C927V997,C927V1095,C927V2079,C927V2175:std_logic_vector(8 downto 0);
signal V542C928,V699C928,V998C928,V1096C928,V2080C928,V2176C928,C928V542,C928V699,C928V998,C928V1096,C928V2080,C928V2176:std_logic_vector(8 downto 0);
signal V543C929,V700C929,V999C929,V1097C929,V2081C929,V2177C929,C929V543,C929V700,C929V999,C929V1097,C929V2081,C929V2177:std_logic_vector(8 downto 0);
signal V544C930,V701C930,V1000C930,V1098C930,V2082C930,V2178C930,C930V544,C930V701,C930V1000,C930V1098,C930V2082,C930V2178:std_logic_vector(8 downto 0);
signal V545C931,V702C931,V1001C931,V1099C931,V2083C931,V2179C931,C931V545,C931V702,C931V1001,C931V1099,C931V2083,C931V2179:std_logic_vector(8 downto 0);
signal V546C932,V703C932,V1002C932,V1100C932,V2084C932,V2180C932,C932V546,C932V703,C932V1002,C932V1100,C932V2084,C932V2180:std_logic_vector(8 downto 0);
signal V547C933,V704C933,V1003C933,V1101C933,V2085C933,V2181C933,C933V547,C933V704,C933V1003,C933V1101,C933V2085,C933V2181:std_logic_vector(8 downto 0);
signal V548C934,V705C934,V1004C934,V1102C934,V2086C934,V2182C934,C934V548,C934V705,C934V1004,C934V1102,C934V2086,C934V2182:std_logic_vector(8 downto 0);
signal V549C935,V706C935,V1005C935,V1103C935,V2087C935,V2183C935,C935V549,C935V706,C935V1005,C935V1103,C935V2087,C935V2183:std_logic_vector(8 downto 0);
signal V550C936,V707C936,V1006C936,V1104C936,V2088C936,V2184C936,C936V550,C936V707,C936V1006,C936V1104,C936V2088,C936V2184:std_logic_vector(8 downto 0);
signal V551C937,V708C937,V1007C937,V1105C937,V2089C937,V2185C937,C937V551,C937V708,C937V1007,C937V1105,C937V2089,C937V2185:std_logic_vector(8 downto 0);
signal V552C938,V709C938,V1008C938,V1106C938,V2090C938,V2186C938,C938V552,C938V709,C938V1008,C938V1106,C938V2090,C938V2186:std_logic_vector(8 downto 0);
signal V553C939,V710C939,V1009C939,V1107C939,V2091C939,V2187C939,C939V553,C939V710,C939V1009,C939V1107,C939V2091,C939V2187:std_logic_vector(8 downto 0);
signal V554C940,V711C940,V1010C940,V1108C940,V2092C940,V2188C940,C940V554,C940V711,C940V1010,C940V1108,C940V2092,C940V2188:std_logic_vector(8 downto 0);
signal V555C941,V712C941,V1011C941,V1109C941,V2093C941,V2189C941,C941V555,C941V712,C941V1011,C941V1109,C941V2093,C941V2189:std_logic_vector(8 downto 0);
signal V556C942,V713C942,V1012C942,V1110C942,V2094C942,V2190C942,C942V556,C942V713,C942V1012,C942V1110,C942V2094,C942V2190:std_logic_vector(8 downto 0);
signal V557C943,V714C943,V1013C943,V1111C943,V2095C943,V2191C943,C943V557,C943V714,C943V1013,C943V1111,C943V2095,C943V2191:std_logic_vector(8 downto 0);
signal V558C944,V715C944,V1014C944,V1112C944,V2096C944,V2192C944,C944V558,C944V715,C944V1014,C944V1112,C944V2096,C944V2192:std_logic_vector(8 downto 0);
signal V559C945,V716C945,V1015C945,V1113C945,V2097C945,V2193C945,C945V559,C945V716,C945V1015,C945V1113,C945V2097,C945V2193:std_logic_vector(8 downto 0);
signal V560C946,V717C946,V1016C946,V1114C946,V2098C946,V2194C946,C946V560,C946V717,C946V1016,C946V1114,C946V2098,C946V2194:std_logic_vector(8 downto 0);
signal V561C947,V718C947,V1017C947,V1115C947,V2099C947,V2195C947,C947V561,C947V718,C947V1017,C947V1115,C947V2099,C947V2195:std_logic_vector(8 downto 0);
signal V562C948,V719C948,V1018C948,V1116C948,V2100C948,V2196C948,C948V562,C948V719,C948V1018,C948V1116,C948V2100,C948V2196:std_logic_vector(8 downto 0);
signal V563C949,V720C949,V1019C949,V1117C949,V2101C949,V2197C949,C949V563,C949V720,C949V1019,C949V1117,C949V2101,C949V2197:std_logic_vector(8 downto 0);
signal V564C950,V721C950,V1020C950,V1118C950,V2102C950,V2198C950,C950V564,C950V721,C950V1020,C950V1118,C950V2102,C950V2198:std_logic_vector(8 downto 0);
signal V565C951,V722C951,V1021C951,V1119C951,V2103C951,V2199C951,C951V565,C951V722,C951V1021,C951V1119,C951V2103,C951V2199:std_logic_vector(8 downto 0);
signal V566C952,V723C952,V1022C952,V1120C952,V2104C952,V2200C952,C952V566,C952V723,C952V1022,C952V1120,C952V2104,C952V2200:std_logic_vector(8 downto 0);
signal V567C953,V724C953,V1023C953,V1121C953,V2105C953,V2201C953,C953V567,C953V724,C953V1023,C953V1121,C953V2105,C953V2201:std_logic_vector(8 downto 0);
signal V568C954,V725C954,V1024C954,V1122C954,V2106C954,V2202C954,C954V568,C954V725,C954V1024,C954V1122,C954V2106,C954V2202:std_logic_vector(8 downto 0);
signal V569C955,V726C955,V1025C955,V1123C955,V2107C955,V2203C955,C955V569,C955V726,C955V1025,C955V1123,C955V2107,C955V2203:std_logic_vector(8 downto 0);
signal V570C956,V727C956,V1026C956,V1124C956,V2108C956,V2204C956,C956V570,C956V727,C956V1026,C956V1124,C956V2108,C956V2204:std_logic_vector(8 downto 0);
signal V571C957,V728C957,V1027C957,V1125C957,V2109C957,V2205C957,C957V571,C957V728,C957V1027,C957V1125,C957V2109,C957V2205:std_logic_vector(8 downto 0);
signal V572C958,V729C958,V1028C958,V1126C958,V2110C958,V2206C958,C958V572,C958V729,C958V1028,C958V1126,C958V2110,C958V2206:std_logic_vector(8 downto 0);
signal V573C959,V730C959,V1029C959,V1127C959,V2111C959,V2207C959,C959V573,C959V730,C959V1029,C959V1127,C959V2111,C959V2207:std_logic_vector(8 downto 0);
signal V574C960,V731C960,V1030C960,V1128C960,V2112C960,V2208C960,C960V574,C960V731,C960V1030,C960V1128,C960V2112,C960V2208:std_logic_vector(8 downto 0);
signal V200C961,V354C961,V808C961,V914C961,V2113C961,V2209C961,C961V200,C961V354,C961V808,C961V914,C961V2113,C961V2209:std_logic_vector(8 downto 0);
signal V201C962,V355C962,V809C962,V915C962,V2114C962,V2210C962,C962V201,C962V355,C962V809,C962V915,C962V2114,C962V2210:std_logic_vector(8 downto 0);
signal V202C963,V356C963,V810C963,V916C963,V2115C963,V2211C963,C963V202,C963V356,C963V810,C963V916,C963V2115,C963V2211:std_logic_vector(8 downto 0);
signal V203C964,V357C964,V811C964,V917C964,V2116C964,V2212C964,C964V203,C964V357,C964V811,C964V917,C964V2116,C964V2212:std_logic_vector(8 downto 0);
signal V204C965,V358C965,V812C965,V918C965,V2117C965,V2213C965,C965V204,C965V358,C965V812,C965V918,C965V2117,C965V2213:std_logic_vector(8 downto 0);
signal V205C966,V359C966,V813C966,V919C966,V2118C966,V2214C966,C966V205,C966V359,C966V813,C966V919,C966V2118,C966V2214:std_logic_vector(8 downto 0);
signal V206C967,V360C967,V814C967,V920C967,V2119C967,V2215C967,C967V206,C967V360,C967V814,C967V920,C967V2119,C967V2215:std_logic_vector(8 downto 0);
signal V207C968,V361C968,V815C968,V921C968,V2120C968,V2216C968,C968V207,C968V361,C968V815,C968V921,C968V2120,C968V2216:std_logic_vector(8 downto 0);
signal V208C969,V362C969,V816C969,V922C969,V2121C969,V2217C969,C969V208,C969V362,C969V816,C969V922,C969V2121,C969V2217:std_logic_vector(8 downto 0);
signal V209C970,V363C970,V817C970,V923C970,V2122C970,V2218C970,C970V209,C970V363,C970V817,C970V923,C970V2122,C970V2218:std_logic_vector(8 downto 0);
signal V210C971,V364C971,V818C971,V924C971,V2123C971,V2219C971,C971V210,C971V364,C971V818,C971V924,C971V2123,C971V2219:std_logic_vector(8 downto 0);
signal V211C972,V365C972,V819C972,V925C972,V2124C972,V2220C972,C972V211,C972V365,C972V819,C972V925,C972V2124,C972V2220:std_logic_vector(8 downto 0);
signal V212C973,V366C973,V820C973,V926C973,V2125C973,V2221C973,C973V212,C973V366,C973V820,C973V926,C973V2125,C973V2221:std_logic_vector(8 downto 0);
signal V213C974,V367C974,V821C974,V927C974,V2126C974,V2222C974,C974V213,C974V367,C974V821,C974V927,C974V2126,C974V2222:std_logic_vector(8 downto 0);
signal V214C975,V368C975,V822C975,V928C975,V2127C975,V2223C975,C975V214,C975V368,C975V822,C975V928,C975V2127,C975V2223:std_logic_vector(8 downto 0);
signal V215C976,V369C976,V823C976,V929C976,V2128C976,V2224C976,C976V215,C976V369,C976V823,C976V929,C976V2128,C976V2224:std_logic_vector(8 downto 0);
signal V216C977,V370C977,V824C977,V930C977,V2129C977,V2225C977,C977V216,C977V370,C977V824,C977V930,C977V2129,C977V2225:std_logic_vector(8 downto 0);
signal V217C978,V371C978,V825C978,V931C978,V2130C978,V2226C978,C978V217,C978V371,C978V825,C978V931,C978V2130,C978V2226:std_logic_vector(8 downto 0);
signal V218C979,V372C979,V826C979,V932C979,V2131C979,V2227C979,C979V218,C979V372,C979V826,C979V932,C979V2131,C979V2227:std_logic_vector(8 downto 0);
signal V219C980,V373C980,V827C980,V933C980,V2132C980,V2228C980,C980V219,C980V373,C980V827,C980V933,C980V2132,C980V2228:std_logic_vector(8 downto 0);
signal V220C981,V374C981,V828C981,V934C981,V2133C981,V2229C981,C981V220,C981V374,C981V828,C981V934,C981V2133,C981V2229:std_logic_vector(8 downto 0);
signal V221C982,V375C982,V829C982,V935C982,V2134C982,V2230C982,C982V221,C982V375,C982V829,C982V935,C982V2134,C982V2230:std_logic_vector(8 downto 0);
signal V222C983,V376C983,V830C983,V936C983,V2135C983,V2231C983,C983V222,C983V376,C983V830,C983V936,C983V2135,C983V2231:std_logic_vector(8 downto 0);
signal V223C984,V377C984,V831C984,V937C984,V2136C984,V2232C984,C984V223,C984V377,C984V831,C984V937,C984V2136,C984V2232:std_logic_vector(8 downto 0);
signal V224C985,V378C985,V832C985,V938C985,V2137C985,V2233C985,C985V224,C985V378,C985V832,C985V938,C985V2137,C985V2233:std_logic_vector(8 downto 0);
signal V225C986,V379C986,V833C986,V939C986,V2138C986,V2234C986,C986V225,C986V379,C986V833,C986V939,C986V2138,C986V2234:std_logic_vector(8 downto 0);
signal V226C987,V380C987,V834C987,V940C987,V2139C987,V2235C987,C987V226,C987V380,C987V834,C987V940,C987V2139,C987V2235:std_logic_vector(8 downto 0);
signal V227C988,V381C988,V835C988,V941C988,V2140C988,V2236C988,C988V227,C988V381,C988V835,C988V941,C988V2140,C988V2236:std_logic_vector(8 downto 0);
signal V228C989,V382C989,V836C989,V942C989,V2141C989,V2237C989,C989V228,C989V382,C989V836,C989V942,C989V2141,C989V2237:std_logic_vector(8 downto 0);
signal V229C990,V383C990,V837C990,V943C990,V2142C990,V2238C990,C990V229,C990V383,C990V837,C990V943,C990V2142,C990V2238:std_logic_vector(8 downto 0);
signal V230C991,V384C991,V838C991,V944C991,V2143C991,V2239C991,C991V230,C991V384,C991V838,C991V944,C991V2143,C991V2239:std_logic_vector(8 downto 0);
signal V231C992,V289C992,V839C992,V945C992,V2144C992,V2240C992,C992V231,C992V289,C992V839,C992V945,C992V2144,C992V2240:std_logic_vector(8 downto 0);
signal V232C993,V290C993,V840C993,V946C993,V2145C993,V2241C993,C993V232,C993V290,C993V840,C993V946,C993V2145,C993V2241:std_logic_vector(8 downto 0);
signal V233C994,V291C994,V841C994,V947C994,V2146C994,V2242C994,C994V233,C994V291,C994V841,C994V947,C994V2146,C994V2242:std_logic_vector(8 downto 0);
signal V234C995,V292C995,V842C995,V948C995,V2147C995,V2243C995,C995V234,C995V292,C995V842,C995V948,C995V2147,C995V2243:std_logic_vector(8 downto 0);
signal V235C996,V293C996,V843C996,V949C996,V2148C996,V2244C996,C996V235,C996V293,C996V843,C996V949,C996V2148,C996V2244:std_logic_vector(8 downto 0);
signal V236C997,V294C997,V844C997,V950C997,V2149C997,V2245C997,C997V236,C997V294,C997V844,C997V950,C997V2149,C997V2245:std_logic_vector(8 downto 0);
signal V237C998,V295C998,V845C998,V951C998,V2150C998,V2246C998,C998V237,C998V295,C998V845,C998V951,C998V2150,C998V2246:std_logic_vector(8 downto 0);
signal V238C999,V296C999,V846C999,V952C999,V2151C999,V2247C999,C999V238,C999V296,C999V846,C999V952,C999V2151,C999V2247:std_logic_vector(8 downto 0);
signal V239C1000,V297C1000,V847C1000,V953C1000,V2152C1000,V2248C1000,C1000V239,C1000V297,C1000V847,C1000V953,C1000V2152,C1000V2248:std_logic_vector(8 downto 0);
signal V240C1001,V298C1001,V848C1001,V954C1001,V2153C1001,V2249C1001,C1001V240,C1001V298,C1001V848,C1001V954,C1001V2153,C1001V2249:std_logic_vector(8 downto 0);
signal V241C1002,V299C1002,V849C1002,V955C1002,V2154C1002,V2250C1002,C1002V241,C1002V299,C1002V849,C1002V955,C1002V2154,C1002V2250:std_logic_vector(8 downto 0);
signal V242C1003,V300C1003,V850C1003,V956C1003,V2155C1003,V2251C1003,C1003V242,C1003V300,C1003V850,C1003V956,C1003V2155,C1003V2251:std_logic_vector(8 downto 0);
signal V243C1004,V301C1004,V851C1004,V957C1004,V2156C1004,V2252C1004,C1004V243,C1004V301,C1004V851,C1004V957,C1004V2156,C1004V2252:std_logic_vector(8 downto 0);
signal V244C1005,V302C1005,V852C1005,V958C1005,V2157C1005,V2253C1005,C1005V244,C1005V302,C1005V852,C1005V958,C1005V2157,C1005V2253:std_logic_vector(8 downto 0);
signal V245C1006,V303C1006,V853C1006,V959C1006,V2158C1006,V2254C1006,C1006V245,C1006V303,C1006V853,C1006V959,C1006V2158,C1006V2254:std_logic_vector(8 downto 0);
signal V246C1007,V304C1007,V854C1007,V960C1007,V2159C1007,V2255C1007,C1007V246,C1007V304,C1007V854,C1007V960,C1007V2159,C1007V2255:std_logic_vector(8 downto 0);
signal V247C1008,V305C1008,V855C1008,V865C1008,V2160C1008,V2256C1008,C1008V247,C1008V305,C1008V855,C1008V865,C1008V2160,C1008V2256:std_logic_vector(8 downto 0);
signal V248C1009,V306C1009,V856C1009,V866C1009,V2161C1009,V2257C1009,C1009V248,C1009V306,C1009V856,C1009V866,C1009V2161,C1009V2257:std_logic_vector(8 downto 0);
signal V249C1010,V307C1010,V857C1010,V867C1010,V2162C1010,V2258C1010,C1010V249,C1010V307,C1010V857,C1010V867,C1010V2162,C1010V2258:std_logic_vector(8 downto 0);
signal V250C1011,V308C1011,V858C1011,V868C1011,V2163C1011,V2259C1011,C1011V250,C1011V308,C1011V858,C1011V868,C1011V2163,C1011V2259:std_logic_vector(8 downto 0);
signal V251C1012,V309C1012,V859C1012,V869C1012,V2164C1012,V2260C1012,C1012V251,C1012V309,C1012V859,C1012V869,C1012V2164,C1012V2260:std_logic_vector(8 downto 0);
signal V252C1013,V310C1013,V860C1013,V870C1013,V2165C1013,V2261C1013,C1013V252,C1013V310,C1013V860,C1013V870,C1013V2165,C1013V2261:std_logic_vector(8 downto 0);
signal V253C1014,V311C1014,V861C1014,V871C1014,V2166C1014,V2262C1014,C1014V253,C1014V311,C1014V861,C1014V871,C1014V2166,C1014V2262:std_logic_vector(8 downto 0);
signal V254C1015,V312C1015,V862C1015,V872C1015,V2167C1015,V2263C1015,C1015V254,C1015V312,C1015V862,C1015V872,C1015V2167,C1015V2263:std_logic_vector(8 downto 0);
signal V255C1016,V313C1016,V863C1016,V873C1016,V2168C1016,V2264C1016,C1016V255,C1016V313,C1016V863,C1016V873,C1016V2168,C1016V2264:std_logic_vector(8 downto 0);
signal V256C1017,V314C1017,V864C1017,V874C1017,V2169C1017,V2265C1017,C1017V256,C1017V314,C1017V864,C1017V874,C1017V2169,C1017V2265:std_logic_vector(8 downto 0);
signal V257C1018,V315C1018,V769C1018,V875C1018,V2170C1018,V2266C1018,C1018V257,C1018V315,C1018V769,C1018V875,C1018V2170,C1018V2266:std_logic_vector(8 downto 0);
signal V258C1019,V316C1019,V770C1019,V876C1019,V2171C1019,V2267C1019,C1019V258,C1019V316,C1019V770,C1019V876,C1019V2171,C1019V2267:std_logic_vector(8 downto 0);
signal V259C1020,V317C1020,V771C1020,V877C1020,V2172C1020,V2268C1020,C1020V259,C1020V317,C1020V771,C1020V877,C1020V2172,C1020V2268:std_logic_vector(8 downto 0);
signal V260C1021,V318C1021,V772C1021,V878C1021,V2173C1021,V2269C1021,C1021V260,C1021V318,C1021V772,C1021V878,C1021V2173,C1021V2269:std_logic_vector(8 downto 0);
signal V261C1022,V319C1022,V773C1022,V879C1022,V2174C1022,V2270C1022,C1022V261,C1022V319,C1022V773,C1022V879,C1022V2174,C1022V2270:std_logic_vector(8 downto 0);
signal V262C1023,V320C1023,V774C1023,V880C1023,V2175C1023,V2271C1023,C1023V262,C1023V320,C1023V774,C1023V880,C1023V2175,C1023V2271:std_logic_vector(8 downto 0);
signal V263C1024,V321C1024,V775C1024,V881C1024,V2176C1024,V2272C1024,C1024V263,C1024V321,C1024V775,C1024V881,C1024V2176,C1024V2272:std_logic_vector(8 downto 0);
signal V264C1025,V322C1025,V776C1025,V882C1025,V2177C1025,V2273C1025,C1025V264,C1025V322,C1025V776,C1025V882,C1025V2177,C1025V2273:std_logic_vector(8 downto 0);
signal V265C1026,V323C1026,V777C1026,V883C1026,V2178C1026,V2274C1026,C1026V265,C1026V323,C1026V777,C1026V883,C1026V2178,C1026V2274:std_logic_vector(8 downto 0);
signal V266C1027,V324C1027,V778C1027,V884C1027,V2179C1027,V2275C1027,C1027V266,C1027V324,C1027V778,C1027V884,C1027V2179,C1027V2275:std_logic_vector(8 downto 0);
signal V267C1028,V325C1028,V779C1028,V885C1028,V2180C1028,V2276C1028,C1028V267,C1028V325,C1028V779,C1028V885,C1028V2180,C1028V2276:std_logic_vector(8 downto 0);
signal V268C1029,V326C1029,V780C1029,V886C1029,V2181C1029,V2277C1029,C1029V268,C1029V326,C1029V780,C1029V886,C1029V2181,C1029V2277:std_logic_vector(8 downto 0);
signal V269C1030,V327C1030,V781C1030,V887C1030,V2182C1030,V2278C1030,C1030V269,C1030V327,C1030V781,C1030V887,C1030V2182,C1030V2278:std_logic_vector(8 downto 0);
signal V270C1031,V328C1031,V782C1031,V888C1031,V2183C1031,V2279C1031,C1031V270,C1031V328,C1031V782,C1031V888,C1031V2183,C1031V2279:std_logic_vector(8 downto 0);
signal V271C1032,V329C1032,V783C1032,V889C1032,V2184C1032,V2280C1032,C1032V271,C1032V329,C1032V783,C1032V889,C1032V2184,C1032V2280:std_logic_vector(8 downto 0);
signal V272C1033,V330C1033,V784C1033,V890C1033,V2185C1033,V2281C1033,C1033V272,C1033V330,C1033V784,C1033V890,C1033V2185,C1033V2281:std_logic_vector(8 downto 0);
signal V273C1034,V331C1034,V785C1034,V891C1034,V2186C1034,V2282C1034,C1034V273,C1034V331,C1034V785,C1034V891,C1034V2186,C1034V2282:std_logic_vector(8 downto 0);
signal V274C1035,V332C1035,V786C1035,V892C1035,V2187C1035,V2283C1035,C1035V274,C1035V332,C1035V786,C1035V892,C1035V2187,C1035V2283:std_logic_vector(8 downto 0);
signal V275C1036,V333C1036,V787C1036,V893C1036,V2188C1036,V2284C1036,C1036V275,C1036V333,C1036V787,C1036V893,C1036V2188,C1036V2284:std_logic_vector(8 downto 0);
signal V276C1037,V334C1037,V788C1037,V894C1037,V2189C1037,V2285C1037,C1037V276,C1037V334,C1037V788,C1037V894,C1037V2189,C1037V2285:std_logic_vector(8 downto 0);
signal V277C1038,V335C1038,V789C1038,V895C1038,V2190C1038,V2286C1038,C1038V277,C1038V335,C1038V789,C1038V895,C1038V2190,C1038V2286:std_logic_vector(8 downto 0);
signal V278C1039,V336C1039,V790C1039,V896C1039,V2191C1039,V2287C1039,C1039V278,C1039V336,C1039V790,C1039V896,C1039V2191,C1039V2287:std_logic_vector(8 downto 0);
signal V279C1040,V337C1040,V791C1040,V897C1040,V2192C1040,V2288C1040,C1040V279,C1040V337,C1040V791,C1040V897,C1040V2192,C1040V2288:std_logic_vector(8 downto 0);
signal V280C1041,V338C1041,V792C1041,V898C1041,V2193C1041,V2289C1041,C1041V280,C1041V338,C1041V792,C1041V898,C1041V2193,C1041V2289:std_logic_vector(8 downto 0);
signal V281C1042,V339C1042,V793C1042,V899C1042,V2194C1042,V2290C1042,C1042V281,C1042V339,C1042V793,C1042V899,C1042V2194,C1042V2290:std_logic_vector(8 downto 0);
signal V282C1043,V340C1043,V794C1043,V900C1043,V2195C1043,V2291C1043,C1043V282,C1043V340,C1043V794,C1043V900,C1043V2195,C1043V2291:std_logic_vector(8 downto 0);
signal V283C1044,V341C1044,V795C1044,V901C1044,V2196C1044,V2292C1044,C1044V283,C1044V341,C1044V795,C1044V901,C1044V2196,C1044V2292:std_logic_vector(8 downto 0);
signal V284C1045,V342C1045,V796C1045,V902C1045,V2197C1045,V2293C1045,C1045V284,C1045V342,C1045V796,C1045V902,C1045V2197,C1045V2293:std_logic_vector(8 downto 0);
signal V285C1046,V343C1046,V797C1046,V903C1046,V2198C1046,V2294C1046,C1046V285,C1046V343,C1046V797,C1046V903,C1046V2198,C1046V2294:std_logic_vector(8 downto 0);
signal V286C1047,V344C1047,V798C1047,V904C1047,V2199C1047,V2295C1047,C1047V286,C1047V344,C1047V798,C1047V904,C1047V2199,C1047V2295:std_logic_vector(8 downto 0);
signal V287C1048,V345C1048,V799C1048,V905C1048,V2200C1048,V2296C1048,C1048V287,C1048V345,C1048V799,C1048V905,C1048V2200,C1048V2296:std_logic_vector(8 downto 0);
signal V288C1049,V346C1049,V800C1049,V906C1049,V2201C1049,V2297C1049,C1049V288,C1049V346,C1049V800,C1049V906,C1049V2201,C1049V2297:std_logic_vector(8 downto 0);
signal V193C1050,V347C1050,V801C1050,V907C1050,V2202C1050,V2298C1050,C1050V193,C1050V347,C1050V801,C1050V907,C1050V2202,C1050V2298:std_logic_vector(8 downto 0);
signal V194C1051,V348C1051,V802C1051,V908C1051,V2203C1051,V2299C1051,C1051V194,C1051V348,C1051V802,C1051V908,C1051V2203,C1051V2299:std_logic_vector(8 downto 0);
signal V195C1052,V349C1052,V803C1052,V909C1052,V2204C1052,V2300C1052,C1052V195,C1052V349,C1052V803,C1052V909,C1052V2204,C1052V2300:std_logic_vector(8 downto 0);
signal V196C1053,V350C1053,V804C1053,V910C1053,V2205C1053,V2301C1053,C1053V196,C1053V350,C1053V804,C1053V910,C1053V2205,C1053V2301:std_logic_vector(8 downto 0);
signal V197C1054,V351C1054,V805C1054,V911C1054,V2206C1054,V2302C1054,C1054V197,C1054V351,C1054V805,C1054V911,C1054V2206,C1054V2302:std_logic_vector(8 downto 0);
signal V198C1055,V352C1055,V806C1055,V912C1055,V2207C1055,V2303C1055,C1055V198,C1055V352,C1055V806,C1055V912,C1055V2207,C1055V2303:std_logic_vector(8 downto 0);
signal V199C1056,V353C1056,V807C1056,V913C1056,V2208C1056,V2304C1056,C1056V199,C1056V353,C1056V807,C1056V913,C1056V2208,C1056V2304:std_logic_vector(8 downto 0);
signal V44C1057,V547C1057,V714C1057,V1083C1057,V1160C1057,V2209C1057,C1057V44,C1057V547,C1057V714,C1057V1083,C1057V1160,C1057V2209:std_logic_vector(8 downto 0);
signal V45C1058,V548C1058,V715C1058,V1084C1058,V1161C1058,V2210C1058,C1058V45,C1058V548,C1058V715,C1058V1084,C1058V1161,C1058V2210:std_logic_vector(8 downto 0);
signal V46C1059,V549C1059,V716C1059,V1085C1059,V1162C1059,V2211C1059,C1059V46,C1059V549,C1059V716,C1059V1085,C1059V1162,C1059V2211:std_logic_vector(8 downto 0);
signal V47C1060,V550C1060,V717C1060,V1086C1060,V1163C1060,V2212C1060,C1060V47,C1060V550,C1060V717,C1060V1086,C1060V1163,C1060V2212:std_logic_vector(8 downto 0);
signal V48C1061,V551C1061,V718C1061,V1087C1061,V1164C1061,V2213C1061,C1061V48,C1061V551,C1061V718,C1061V1087,C1061V1164,C1061V2213:std_logic_vector(8 downto 0);
signal V49C1062,V552C1062,V719C1062,V1088C1062,V1165C1062,V2214C1062,C1062V49,C1062V552,C1062V719,C1062V1088,C1062V1165,C1062V2214:std_logic_vector(8 downto 0);
signal V50C1063,V553C1063,V720C1063,V1089C1063,V1166C1063,V2215C1063,C1063V50,C1063V553,C1063V720,C1063V1089,C1063V1166,C1063V2215:std_logic_vector(8 downto 0);
signal V51C1064,V554C1064,V721C1064,V1090C1064,V1167C1064,V2216C1064,C1064V51,C1064V554,C1064V721,C1064V1090,C1064V1167,C1064V2216:std_logic_vector(8 downto 0);
signal V52C1065,V555C1065,V722C1065,V1091C1065,V1168C1065,V2217C1065,C1065V52,C1065V555,C1065V722,C1065V1091,C1065V1168,C1065V2217:std_logic_vector(8 downto 0);
signal V53C1066,V556C1066,V723C1066,V1092C1066,V1169C1066,V2218C1066,C1066V53,C1066V556,C1066V723,C1066V1092,C1066V1169,C1066V2218:std_logic_vector(8 downto 0);
signal V54C1067,V557C1067,V724C1067,V1093C1067,V1170C1067,V2219C1067,C1067V54,C1067V557,C1067V724,C1067V1093,C1067V1170,C1067V2219:std_logic_vector(8 downto 0);
signal V55C1068,V558C1068,V725C1068,V1094C1068,V1171C1068,V2220C1068,C1068V55,C1068V558,C1068V725,C1068V1094,C1068V1171,C1068V2220:std_logic_vector(8 downto 0);
signal V56C1069,V559C1069,V726C1069,V1095C1069,V1172C1069,V2221C1069,C1069V56,C1069V559,C1069V726,C1069V1095,C1069V1172,C1069V2221:std_logic_vector(8 downto 0);
signal V57C1070,V560C1070,V727C1070,V1096C1070,V1173C1070,V2222C1070,C1070V57,C1070V560,C1070V727,C1070V1096,C1070V1173,C1070V2222:std_logic_vector(8 downto 0);
signal V58C1071,V561C1071,V728C1071,V1097C1071,V1174C1071,V2223C1071,C1071V58,C1071V561,C1071V728,C1071V1097,C1071V1174,C1071V2223:std_logic_vector(8 downto 0);
signal V59C1072,V562C1072,V729C1072,V1098C1072,V1175C1072,V2224C1072,C1072V59,C1072V562,C1072V729,C1072V1098,C1072V1175,C1072V2224:std_logic_vector(8 downto 0);
signal V60C1073,V563C1073,V730C1073,V1099C1073,V1176C1073,V2225C1073,C1073V60,C1073V563,C1073V730,C1073V1099,C1073V1176,C1073V2225:std_logic_vector(8 downto 0);
signal V61C1074,V564C1074,V731C1074,V1100C1074,V1177C1074,V2226C1074,C1074V61,C1074V564,C1074V731,C1074V1100,C1074V1177,C1074V2226:std_logic_vector(8 downto 0);
signal V62C1075,V565C1075,V732C1075,V1101C1075,V1178C1075,V2227C1075,C1075V62,C1075V565,C1075V732,C1075V1101,C1075V1178,C1075V2227:std_logic_vector(8 downto 0);
signal V63C1076,V566C1076,V733C1076,V1102C1076,V1179C1076,V2228C1076,C1076V63,C1076V566,C1076V733,C1076V1102,C1076V1179,C1076V2228:std_logic_vector(8 downto 0);
signal V64C1077,V567C1077,V734C1077,V1103C1077,V1180C1077,V2229C1077,C1077V64,C1077V567,C1077V734,C1077V1103,C1077V1180,C1077V2229:std_logic_vector(8 downto 0);
signal V65C1078,V568C1078,V735C1078,V1104C1078,V1181C1078,V2230C1078,C1078V65,C1078V568,C1078V735,C1078V1104,C1078V1181,C1078V2230:std_logic_vector(8 downto 0);
signal V66C1079,V569C1079,V736C1079,V1105C1079,V1182C1079,V2231C1079,C1079V66,C1079V569,C1079V736,C1079V1105,C1079V1182,C1079V2231:std_logic_vector(8 downto 0);
signal V67C1080,V570C1080,V737C1080,V1106C1080,V1183C1080,V2232C1080,C1080V67,C1080V570,C1080V737,C1080V1106,C1080V1183,C1080V2232:std_logic_vector(8 downto 0);
signal V68C1081,V571C1081,V738C1081,V1107C1081,V1184C1081,V2233C1081,C1081V68,C1081V571,C1081V738,C1081V1107,C1081V1184,C1081V2233:std_logic_vector(8 downto 0);
signal V69C1082,V572C1082,V739C1082,V1108C1082,V1185C1082,V2234C1082,C1082V69,C1082V572,C1082V739,C1082V1108,C1082V1185,C1082V2234:std_logic_vector(8 downto 0);
signal V70C1083,V573C1083,V740C1083,V1109C1083,V1186C1083,V2235C1083,C1083V70,C1083V573,C1083V740,C1083V1109,C1083V1186,C1083V2235:std_logic_vector(8 downto 0);
signal V71C1084,V574C1084,V741C1084,V1110C1084,V1187C1084,V2236C1084,C1084V71,C1084V574,C1084V741,C1084V1110,C1084V1187,C1084V2236:std_logic_vector(8 downto 0);
signal V72C1085,V575C1085,V742C1085,V1111C1085,V1188C1085,V2237C1085,C1085V72,C1085V575,C1085V742,C1085V1111,C1085V1188,C1085V2237:std_logic_vector(8 downto 0);
signal V73C1086,V576C1086,V743C1086,V1112C1086,V1189C1086,V2238C1086,C1086V73,C1086V576,C1086V743,C1086V1112,C1086V1189,C1086V2238:std_logic_vector(8 downto 0);
signal V74C1087,V481C1087,V744C1087,V1113C1087,V1190C1087,V2239C1087,C1087V74,C1087V481,C1087V744,C1087V1113,C1087V1190,C1087V2239:std_logic_vector(8 downto 0);
signal V75C1088,V482C1088,V745C1088,V1114C1088,V1191C1088,V2240C1088,C1088V75,C1088V482,C1088V745,C1088V1114,C1088V1191,C1088V2240:std_logic_vector(8 downto 0);
signal V76C1089,V483C1089,V746C1089,V1115C1089,V1192C1089,V2241C1089,C1089V76,C1089V483,C1089V746,C1089V1115,C1089V1192,C1089V2241:std_logic_vector(8 downto 0);
signal V77C1090,V484C1090,V747C1090,V1116C1090,V1193C1090,V2242C1090,C1090V77,C1090V484,C1090V747,C1090V1116,C1090V1193,C1090V2242:std_logic_vector(8 downto 0);
signal V78C1091,V485C1091,V748C1091,V1117C1091,V1194C1091,V2243C1091,C1091V78,C1091V485,C1091V748,C1091V1117,C1091V1194,C1091V2243:std_logic_vector(8 downto 0);
signal V79C1092,V486C1092,V749C1092,V1118C1092,V1195C1092,V2244C1092,C1092V79,C1092V486,C1092V749,C1092V1118,C1092V1195,C1092V2244:std_logic_vector(8 downto 0);
signal V80C1093,V487C1093,V750C1093,V1119C1093,V1196C1093,V2245C1093,C1093V80,C1093V487,C1093V750,C1093V1119,C1093V1196,C1093V2245:std_logic_vector(8 downto 0);
signal V81C1094,V488C1094,V751C1094,V1120C1094,V1197C1094,V2246C1094,C1094V81,C1094V488,C1094V751,C1094V1120,C1094V1197,C1094V2246:std_logic_vector(8 downto 0);
signal V82C1095,V489C1095,V752C1095,V1121C1095,V1198C1095,V2247C1095,C1095V82,C1095V489,C1095V752,C1095V1121,C1095V1198,C1095V2247:std_logic_vector(8 downto 0);
signal V83C1096,V490C1096,V753C1096,V1122C1096,V1199C1096,V2248C1096,C1096V83,C1096V490,C1096V753,C1096V1122,C1096V1199,C1096V2248:std_logic_vector(8 downto 0);
signal V84C1097,V491C1097,V754C1097,V1123C1097,V1200C1097,V2249C1097,C1097V84,C1097V491,C1097V754,C1097V1123,C1097V1200,C1097V2249:std_logic_vector(8 downto 0);
signal V85C1098,V492C1098,V755C1098,V1124C1098,V1201C1098,V2250C1098,C1098V85,C1098V492,C1098V755,C1098V1124,C1098V1201,C1098V2250:std_logic_vector(8 downto 0);
signal V86C1099,V493C1099,V756C1099,V1125C1099,V1202C1099,V2251C1099,C1099V86,C1099V493,C1099V756,C1099V1125,C1099V1202,C1099V2251:std_logic_vector(8 downto 0);
signal V87C1100,V494C1100,V757C1100,V1126C1100,V1203C1100,V2252C1100,C1100V87,C1100V494,C1100V757,C1100V1126,C1100V1203,C1100V2252:std_logic_vector(8 downto 0);
signal V88C1101,V495C1101,V758C1101,V1127C1101,V1204C1101,V2253C1101,C1101V88,C1101V495,C1101V758,C1101V1127,C1101V1204,C1101V2253:std_logic_vector(8 downto 0);
signal V89C1102,V496C1102,V759C1102,V1128C1102,V1205C1102,V2254C1102,C1102V89,C1102V496,C1102V759,C1102V1128,C1102V1205,C1102V2254:std_logic_vector(8 downto 0);
signal V90C1103,V497C1103,V760C1103,V1129C1103,V1206C1103,V2255C1103,C1103V90,C1103V497,C1103V760,C1103V1129,C1103V1206,C1103V2255:std_logic_vector(8 downto 0);
signal V91C1104,V498C1104,V761C1104,V1130C1104,V1207C1104,V2256C1104,C1104V91,C1104V498,C1104V761,C1104V1130,C1104V1207,C1104V2256:std_logic_vector(8 downto 0);
signal V92C1105,V499C1105,V762C1105,V1131C1105,V1208C1105,V2257C1105,C1105V92,C1105V499,C1105V762,C1105V1131,C1105V1208,C1105V2257:std_logic_vector(8 downto 0);
signal V93C1106,V500C1106,V763C1106,V1132C1106,V1209C1106,V2258C1106,C1106V93,C1106V500,C1106V763,C1106V1132,C1106V1209,C1106V2258:std_logic_vector(8 downto 0);
signal V94C1107,V501C1107,V764C1107,V1133C1107,V1210C1107,V2259C1107,C1107V94,C1107V501,C1107V764,C1107V1133,C1107V1210,C1107V2259:std_logic_vector(8 downto 0);
signal V95C1108,V502C1108,V765C1108,V1134C1108,V1211C1108,V2260C1108,C1108V95,C1108V502,C1108V765,C1108V1134,C1108V1211,C1108V2260:std_logic_vector(8 downto 0);
signal V96C1109,V503C1109,V766C1109,V1135C1109,V1212C1109,V2261C1109,C1109V96,C1109V503,C1109V766,C1109V1135,C1109V1212,C1109V2261:std_logic_vector(8 downto 0);
signal V1C1110,V504C1110,V767C1110,V1136C1110,V1213C1110,V2262C1110,C1110V1,C1110V504,C1110V767,C1110V1136,C1110V1213,C1110V2262:std_logic_vector(8 downto 0);
signal V2C1111,V505C1111,V768C1111,V1137C1111,V1214C1111,V2263C1111,C1111V2,C1111V505,C1111V768,C1111V1137,C1111V1214,C1111V2263:std_logic_vector(8 downto 0);
signal V3C1112,V506C1112,V673C1112,V1138C1112,V1215C1112,V2264C1112,C1112V3,C1112V506,C1112V673,C1112V1138,C1112V1215,C1112V2264:std_logic_vector(8 downto 0);
signal V4C1113,V507C1113,V674C1113,V1139C1113,V1216C1113,V2265C1113,C1113V4,C1113V507,C1113V674,C1113V1139,C1113V1216,C1113V2265:std_logic_vector(8 downto 0);
signal V5C1114,V508C1114,V675C1114,V1140C1114,V1217C1114,V2266C1114,C1114V5,C1114V508,C1114V675,C1114V1140,C1114V1217,C1114V2266:std_logic_vector(8 downto 0);
signal V6C1115,V509C1115,V676C1115,V1141C1115,V1218C1115,V2267C1115,C1115V6,C1115V509,C1115V676,C1115V1141,C1115V1218,C1115V2267:std_logic_vector(8 downto 0);
signal V7C1116,V510C1116,V677C1116,V1142C1116,V1219C1116,V2268C1116,C1116V7,C1116V510,C1116V677,C1116V1142,C1116V1219,C1116V2268:std_logic_vector(8 downto 0);
signal V8C1117,V511C1117,V678C1117,V1143C1117,V1220C1117,V2269C1117,C1117V8,C1117V511,C1117V678,C1117V1143,C1117V1220,C1117V2269:std_logic_vector(8 downto 0);
signal V9C1118,V512C1118,V679C1118,V1144C1118,V1221C1118,V2270C1118,C1118V9,C1118V512,C1118V679,C1118V1144,C1118V1221,C1118V2270:std_logic_vector(8 downto 0);
signal V10C1119,V513C1119,V680C1119,V1145C1119,V1222C1119,V2271C1119,C1119V10,C1119V513,C1119V680,C1119V1145,C1119V1222,C1119V2271:std_logic_vector(8 downto 0);
signal V11C1120,V514C1120,V681C1120,V1146C1120,V1223C1120,V2272C1120,C1120V11,C1120V514,C1120V681,C1120V1146,C1120V1223,C1120V2272:std_logic_vector(8 downto 0);
signal V12C1121,V515C1121,V682C1121,V1147C1121,V1224C1121,V2273C1121,C1121V12,C1121V515,C1121V682,C1121V1147,C1121V1224,C1121V2273:std_logic_vector(8 downto 0);
signal V13C1122,V516C1122,V683C1122,V1148C1122,V1225C1122,V2274C1122,C1122V13,C1122V516,C1122V683,C1122V1148,C1122V1225,C1122V2274:std_logic_vector(8 downto 0);
signal V14C1123,V517C1123,V684C1123,V1149C1123,V1226C1123,V2275C1123,C1123V14,C1123V517,C1123V684,C1123V1149,C1123V1226,C1123V2275:std_logic_vector(8 downto 0);
signal V15C1124,V518C1124,V685C1124,V1150C1124,V1227C1124,V2276C1124,C1124V15,C1124V518,C1124V685,C1124V1150,C1124V1227,C1124V2276:std_logic_vector(8 downto 0);
signal V16C1125,V519C1125,V686C1125,V1151C1125,V1228C1125,V2277C1125,C1125V16,C1125V519,C1125V686,C1125V1151,C1125V1228,C1125V2277:std_logic_vector(8 downto 0);
signal V17C1126,V520C1126,V687C1126,V1152C1126,V1229C1126,V2278C1126,C1126V17,C1126V520,C1126V687,C1126V1152,C1126V1229,C1126V2278:std_logic_vector(8 downto 0);
signal V18C1127,V521C1127,V688C1127,V1057C1127,V1230C1127,V2279C1127,C1127V18,C1127V521,C1127V688,C1127V1057,C1127V1230,C1127V2279:std_logic_vector(8 downto 0);
signal V19C1128,V522C1128,V689C1128,V1058C1128,V1231C1128,V2280C1128,C1128V19,C1128V522,C1128V689,C1128V1058,C1128V1231,C1128V2280:std_logic_vector(8 downto 0);
signal V20C1129,V523C1129,V690C1129,V1059C1129,V1232C1129,V2281C1129,C1129V20,C1129V523,C1129V690,C1129V1059,C1129V1232,C1129V2281:std_logic_vector(8 downto 0);
signal V21C1130,V524C1130,V691C1130,V1060C1130,V1233C1130,V2282C1130,C1130V21,C1130V524,C1130V691,C1130V1060,C1130V1233,C1130V2282:std_logic_vector(8 downto 0);
signal V22C1131,V525C1131,V692C1131,V1061C1131,V1234C1131,V2283C1131,C1131V22,C1131V525,C1131V692,C1131V1061,C1131V1234,C1131V2283:std_logic_vector(8 downto 0);
signal V23C1132,V526C1132,V693C1132,V1062C1132,V1235C1132,V2284C1132,C1132V23,C1132V526,C1132V693,C1132V1062,C1132V1235,C1132V2284:std_logic_vector(8 downto 0);
signal V24C1133,V527C1133,V694C1133,V1063C1133,V1236C1133,V2285C1133,C1133V24,C1133V527,C1133V694,C1133V1063,C1133V1236,C1133V2285:std_logic_vector(8 downto 0);
signal V25C1134,V528C1134,V695C1134,V1064C1134,V1237C1134,V2286C1134,C1134V25,C1134V528,C1134V695,C1134V1064,C1134V1237,C1134V2286:std_logic_vector(8 downto 0);
signal V26C1135,V529C1135,V696C1135,V1065C1135,V1238C1135,V2287C1135,C1135V26,C1135V529,C1135V696,C1135V1065,C1135V1238,C1135V2287:std_logic_vector(8 downto 0);
signal V27C1136,V530C1136,V697C1136,V1066C1136,V1239C1136,V2288C1136,C1136V27,C1136V530,C1136V697,C1136V1066,C1136V1239,C1136V2288:std_logic_vector(8 downto 0);
signal V28C1137,V531C1137,V698C1137,V1067C1137,V1240C1137,V2289C1137,C1137V28,C1137V531,C1137V698,C1137V1067,C1137V1240,C1137V2289:std_logic_vector(8 downto 0);
signal V29C1138,V532C1138,V699C1138,V1068C1138,V1241C1138,V2290C1138,C1138V29,C1138V532,C1138V699,C1138V1068,C1138V1241,C1138V2290:std_logic_vector(8 downto 0);
signal V30C1139,V533C1139,V700C1139,V1069C1139,V1242C1139,V2291C1139,C1139V30,C1139V533,C1139V700,C1139V1069,C1139V1242,C1139V2291:std_logic_vector(8 downto 0);
signal V31C1140,V534C1140,V701C1140,V1070C1140,V1243C1140,V2292C1140,C1140V31,C1140V534,C1140V701,C1140V1070,C1140V1243,C1140V2292:std_logic_vector(8 downto 0);
signal V32C1141,V535C1141,V702C1141,V1071C1141,V1244C1141,V2293C1141,C1141V32,C1141V535,C1141V702,C1141V1071,C1141V1244,C1141V2293:std_logic_vector(8 downto 0);
signal V33C1142,V536C1142,V703C1142,V1072C1142,V1245C1142,V2294C1142,C1142V33,C1142V536,C1142V703,C1142V1072,C1142V1245,C1142V2294:std_logic_vector(8 downto 0);
signal V34C1143,V537C1143,V704C1143,V1073C1143,V1246C1143,V2295C1143,C1143V34,C1143V537,C1143V704,C1143V1073,C1143V1246,C1143V2295:std_logic_vector(8 downto 0);
signal V35C1144,V538C1144,V705C1144,V1074C1144,V1247C1144,V2296C1144,C1144V35,C1144V538,C1144V705,C1144V1074,C1144V1247,C1144V2296:std_logic_vector(8 downto 0);
signal V36C1145,V539C1145,V706C1145,V1075C1145,V1248C1145,V2297C1145,C1145V36,C1145V539,C1145V706,C1145V1075,C1145V1248,C1145V2297:std_logic_vector(8 downto 0);
signal V37C1146,V540C1146,V707C1146,V1076C1146,V1153C1146,V2298C1146,C1146V37,C1146V540,C1146V707,C1146V1076,C1146V1153,C1146V2298:std_logic_vector(8 downto 0);
signal V38C1147,V541C1147,V708C1147,V1077C1147,V1154C1147,V2299C1147,C1147V38,C1147V541,C1147V708,C1147V1077,C1147V1154,C1147V2299:std_logic_vector(8 downto 0);
signal V39C1148,V542C1148,V709C1148,V1078C1148,V1155C1148,V2300C1148,C1148V39,C1148V542,C1148V709,C1148V1078,C1148V1155,C1148V2300:std_logic_vector(8 downto 0);
signal V40C1149,V543C1149,V710C1149,V1079C1149,V1156C1149,V2301C1149,C1149V40,C1149V543,C1149V710,C1149V1079,C1149V1156,C1149V2301:std_logic_vector(8 downto 0);
signal V41C1150,V544C1150,V711C1150,V1080C1150,V1157C1150,V2302C1150,C1150V41,C1150V544,C1150V711,C1150V1080,C1150V1157,C1150V2302:std_logic_vector(8 downto 0);
signal V42C1151,V545C1151,V712C1151,V1081C1151,V1158C1151,V2303C1151,C1151V42,C1151V545,C1151V712,C1151V1081,C1151V1158,C1151V2303:std_logic_vector(8 downto 0);
signal V43C1152,V546C1152,V713C1152,V1082C1152,V1159C1152,V2304C1152,C1152V43,C1152V546,C1152V713,C1152V1082,C1152V1159,C1152V2304:std_logic_vector(8 downto 0);
signal SI1,SI2,SI3,SI4,SI5,SI6,SI7,SI8,SI9,SI10,SI11,SI12,SI13,SI14,SI15,SI16,SI17,SI18,SI19,SI20,SI21,SI22,SI23,SI24,SI25,SI26,SI27,SI28,SI29,SI30,SI31,SI32,SI33,SI34,SI35,SI36,SI37,SI38,SI39,SI40,SI41,SI42,SI43,SI44,SI45,SI46,SI47,SI48,SI49,SI50,SI51,SI52,SI53,SI54,SI55,SI56,SI57,SI58,SI59,SI60,SI61,SI62,SI63,SI64,SI65,SI66,SI67,SI68,SI69,SI70,SI71,SI72,SI73,SI74,SI75,SI76,SI77,SI78,SI79,SI80,SI81,SI82,SI83,SI84,SI85,SI86,SI87,SI88,SI89,SI90,SI91,SI92,SI93,SI94,SI95,SI96,SI97,SI98,SI99,SI100,SI101,SI102,SI103,SI104,SI105,SI106,SI107,SI108,SI109,SI110,SI111,SI112,SI113,SI114,SI115,SI116,SI117,SI118,SI119,SI120,SI121,SI122,SI123,SI124,SI125,SI126,SI127,SI128,SI129,SI130,SI131,SI132,SI133,SI134,SI135,SI136,SI137,SI138,SI139,SI140,SI141,SI142,SI143,SI144,SI145,SI146,SI147,SI148,SI149,SI150,SI151,SI152,SI153,SI154,SI155,SI156,SI157,SI158,SI159,SI160,SI161,SI162,SI163,SI164,SI165,SI166,SI167,SI168,SI169,SI170,SI171,SI172,SI173,SI174,SI175,SI176,SI177,SI178,SI179,SI180,SI181,SI182,SI183,SI184,SI185,SI186,SI187,SI188,SI189,SI190,SI191,SI192,SI193,SI194,SI195,SI196,SI197,SI198,SI199,SI200,SI201,SI202,SI203,SI204,SI205,SI206,SI207,SI208,SI209,SI210,SI211,SI212,SI213,SI214,SI215,SI216,SI217,SI218,SI219,SI220,SI221,SI222,SI223,SI224,SI225,SI226,SI227,SI228,SI229,SI230,SI231,SI232,SI233,SI234,SI235,SI236,SI237,SI238,SI239,SI240,SI241,SI242,SI243,SI244,SI245,SI246,SI247,SI248,SI249,SI250,SI251,SI252,SI253,SI254,SI255,SI256,SI257,SI258,SI259,SI260,SI261,SI262,SI263,SI264,SI265,SI266,SI267,SI268,SI269,SI270,SI271,SI272,SI273,SI274,SI275,SI276,SI277,SI278,SI279,SI280,SI281,SI282,SI283,SI284,SI285,SI286,SI287,SI288,SI289,SI290,SI291,SI292,SI293,SI294,SI295,SI296,SI297,SI298,SI299,SI300,SI301,SI302,SI303,SI304,SI305,SI306,SI307,SI308,SI309,SI310,SI311,SI312,SI313,SI314,SI315,SI316,SI317,SI318,SI319,SI320,SI321,SI322,SI323,SI324,SI325,SI326,SI327,SI328,SI329,SI330,SI331,SI332,SI333,SI334,SI335,SI336,SI337,SI338,SI339,SI340,SI341,SI342,SI343,SI344,SI345,SI346,SI347,SI348,SI349,SI350,SI351,SI352,SI353,SI354,SI355,SI356,SI357,SI358,SI359,SI360,SI361,SI362,SI363,SI364,SI365,SI366,SI367,SI368,SI369,SI370,SI371,SI372,SI373,SI374,SI375,SI376,SI377,SI378,SI379,SI380,SI381,SI382,SI383,SI384,SI385,SI386,SI387,SI388,SI389,SI390,SI391,SI392,SI393,SI394,SI395,SI396,SI397,SI398,SI399,SI400,SI401,SI402,SI403,SI404,SI405,SI406,SI407,SI408,SI409,SI410,SI411,SI412,SI413,SI414,SI415,SI416,SI417,SI418,SI419,SI420,SI421,SI422,SI423,SI424,SI425,SI426,SI427,SI428,SI429,SI430,SI431,SI432,SI433,SI434,SI435,SI436,SI437,SI438,SI439,SI440,SI441,SI442,SI443,SI444,SI445,SI446,SI447,SI448,SI449,SI450,SI451,SI452,SI453,SI454,SI455,SI456,SI457,SI458,SI459,SI460,SI461,SI462,SI463,SI464,SI465,SI466,SI467,SI468,SI469,SI470,SI471,SI472,SI473,SI474,SI475,SI476,SI477,SI478,SI479,SI480,SI481,SI482,SI483,SI484,SI485,SI486,SI487,SI488,SI489,SI490,SI491,SI492,SI493,SI494,SI495,SI496,SI497,SI498,SI499,SI500,SI501,SI502,SI503,SI504,SI505,SI506,SI507,SI508,SI509,SI510,SI511,SI512,SI513,SI514,SI515,SI516,SI517,SI518,SI519,SI520,SI521,SI522,SI523,SI524,SI525,SI526,SI527,SI528,SI529,SI530,SI531,SI532,SI533,SI534,SI535,SI536,SI537,SI538,SI539,SI540,SI541,SI542,SI543,SI544,SI545,SI546,SI547,SI548,SI549,SI550,SI551,SI552,SI553,SI554,SI555,SI556,SI557,SI558,SI559,SI560,SI561,SI562,SI563,SI564,SI565,SI566,SI567,SI568,SI569,SI570,SI571,SI572,SI573,SI574,SI575,SI576,SI577,SI578,SI579,SI580,SI581,SI582,SI583,SI584,SI585,SI586,SI587,SI588,SI589,SI590,SI591,SI592,SI593,SI594,SI595,SI596,SI597,SI598,SI599,SI600,SI601,SI602,SI603,SI604,SI605,SI606,SI607,SI608,SI609,SI610,SI611,SI612,SI613,SI614,SI615,SI616,SI617,SI618,SI619,SI620,SI621,SI622,SI623,SI624,SI625,SI626,SI627,SI628,SI629,SI630,SI631,SI632,SI633,SI634,SI635,SI636,SI637,SI638,SI639,SI640,SI641,SI642,SI643,SI644,SI645,SI646,SI647,SI648,SI649,SI650,SI651,SI652,SI653,SI654,SI655,SI656,SI657,SI658,SI659,SI660,SI661,SI662,SI663,SI664,SI665,SI666,SI667,SI668,SI669,SI670,SI671,SI672,SI673,SI674,SI675,SI676,SI677,SI678,SI679,SI680,SI681,SI682,SI683,SI684,SI685,SI686,SI687,SI688,SI689,SI690,SI691,SI692,SI693,SI694,SI695,SI696,SI697,SI698,SI699,SI700,SI701,SI702,SI703,SI704,SI705,SI706,SI707,SI708,SI709,SI710,SI711,SI712,SI713,SI714,SI715,SI716,SI717,SI718,SI719,SI720,SI721,SI722,SI723,SI724,SI725,SI726,SI727,SI728,SI729,SI730,SI731,SI732,SI733,SI734,SI735,SI736,SI737,SI738,SI739,SI740,SI741,SI742,SI743,SI744,SI745,SI746,SI747,SI748,SI749,SI750,SI751,SI752,SI753,SI754,SI755,SI756,SI757,SI758,SI759,SI760,SI761,SI762,SI763,SI764,SI765,SI766,SI767,SI768,SI769,SI770,SI771,SI772,SI773,SI774,SI775,SI776,SI777,SI778,SI779,SI780,SI781,SI782,SI783,SI784,SI785,SI786,SI787,SI788,SI789,SI790,SI791,SI792,SI793,SI794,SI795,SI796,SI797,SI798,SI799,SI800,SI801,SI802,SI803,SI804,SI805,SI806,SI807,SI808,SI809,SI810,SI811,SI812,SI813,SI814,SI815,SI816,SI817,SI818,SI819,SI820,SI821,SI822,SI823,SI824,SI825,SI826,SI827,SI828,SI829,SI830,SI831,SI832,SI833,SI834,SI835,SI836,SI837,SI838,SI839,SI840,SI841,SI842,SI843,SI844,SI845,SI846,SI847,SI848,SI849,SI850,SI851,SI852,SI853,SI854,SI855,SI856,SI857,SI858,SI859,SI860,SI861,SI862,SI863,SI864,SI865,SI866,SI867,SI868,SI869,SI870,SI871,SI872,SI873,SI874,SI875,SI876,SI877,SI878,SI879,SI880,SI881,SI882,SI883,SI884,SI885,SI886,SI887,SI888,SI889,SI890,SI891,SI892,SI893,SI894,SI895,SI896,SI897,SI898,SI899,SI900,SI901,SI902,SI903,SI904,SI905,SI906,SI907,SI908,SI909,SI910,SI911,SI912,SI913,SI914,SI915,SI916,SI917,SI918,SI919,SI920,SI921,SI922,SI923,SI924,SI925,SI926,SI927,SI928,SI929,SI930,SI931,SI932,SI933,SI934,SI935,SI936,SI937,SI938,SI939,SI940,SI941,SI942,SI943,SI944,SI945,SI946,SI947,SI948,SI949,SI950,SI951,SI952,SI953,SI954,SI955,SI956,SI957,SI958,SI959,SI960,SI961,SI962,SI963,SI964,SI965,SI966,SI967,SI968,SI969,SI970,SI971,SI972,SI973,SI974,SI975,SI976,SI977,SI978,SI979,SI980,SI981,SI982,SI983,SI984,SI985,SI986,SI987,SI988,SI989,SI990,SI991,SI992,SI993,SI994,SI995,SI996,SI997,SI998,SI999,SI1000,SI1001,SI1002,SI1003,SI1004,SI1005,SI1006,SI1007,SI1008,SI1009,SI1010,SI1011,SI1012,SI1013,SI1014,SI1015,SI1016,SI1017,SI1018,SI1019,SI1020,SI1021,SI1022,SI1023,SI1024,SI1025,SI1026,SI1027,SI1028,SI1029,SI1030,SI1031,SI1032,SI1033,SI1034,SI1035,SI1036,SI1037,SI1038,SI1039,SI1040,SI1041,SI1042,SI1043,SI1044,SI1045,SI1046,SI1047,SI1048,SI1049,SI1050,SI1051,SI1052,SI1053,SI1054,SI1055,SI1056,SI1057,SI1058,SI1059,SI1060,SI1061,SI1062,SI1063,SI1064,SI1065,SI1066,SI1067,SI1068,SI1069,SI1070,SI1071,SI1072,SI1073,SI1074,SI1075,SI1076,SI1077,SI1078,SI1079,SI1080,SI1081,SI1082,SI1083,SI1084,SI1085,SI1086,SI1087,SI1088,SI1089,SI1090,SI1091,SI1092,SI1093,SI1094,SI1095,SI1096,SI1097,SI1098,SI1099,SI1100,SI1101,SI1102,SI1103,SI1104,SI1105,SI1106,SI1107,SI1108,SI1109,SI1110,SI1111,SI1112,SI1113,SI1114,SI1115,SI1116,SI1117,SI1118,SI1119,SI1120,SI1121,SI1122,SI1123,SI1124,SI1125,SI1126,SI1127,SI1128,SI1129,SI1130,SI1131,SI1132,SI1133,SI1134,SI1135,SI1136,SI1137,SI1138,SI1139,SI1140,SI1141,SI1142,SI1143,SI1144,SI1145,SI1146,SI1147,SI1148,SI1149,SI1150,SI1151,SI1152,SI1153,SI1154,SI1155,SI1156,SI1157,SI1158,SI1159,SI1160,SI1161,SI1162,SI1163,SI1164,SI1165,SI1166,SI1167,SI1168,SI1169,SI1170,SI1171,SI1172,SI1173,SI1174,SI1175,SI1176,SI1177,SI1178,SI1179,SI1180,SI1181,SI1182,SI1183,SI1184,SI1185,SI1186,SI1187,SI1188,SI1189,SI1190,SI1191,SI1192,SI1193,SI1194,SI1195,SI1196,SI1197,SI1198,SI1199,SI1200,SI1201,SI1202,SI1203,SI1204,SI1205,SI1206,SI1207,SI1208,SI1209,SI1210,SI1211,SI1212,SI1213,SI1214,SI1215,SI1216,SI1217,SI1218,SI1219,SI1220,SI1221,SI1222,SI1223,SI1224,SI1225,SI1226,SI1227,SI1228,SI1229,SI1230,SI1231,SI1232,SI1233,SI1234,SI1235,SI1236,SI1237,SI1238,SI1239,SI1240,SI1241,SI1242,SI1243,SI1244,SI1245,SI1246,SI1247,SI1248,SI1249,SI1250,SI1251,SI1252,SI1253,SI1254,SI1255,SI1256,SI1257,SI1258,SI1259,SI1260,SI1261,SI1262,SI1263,SI1264,SI1265,SI1266,SI1267,SI1268,SI1269,SI1270,SI1271,SI1272,SI1273,SI1274,SI1275,SI1276,SI1277,SI1278,SI1279,SI1280,SI1281,SI1282,SI1283,SI1284,SI1285,SI1286,SI1287,SI1288,SI1289,SI1290,SI1291,SI1292,SI1293,SI1294,SI1295,SI1296,SI1297,SI1298,SI1299,SI1300,SI1301,SI1302,SI1303,SI1304,SI1305,SI1306,SI1307,SI1308,SI1309,SI1310,SI1311,SI1312,SI1313,SI1314,SI1315,SI1316,SI1317,SI1318,SI1319,SI1320,SI1321,SI1322,SI1323,SI1324,SI1325,SI1326,SI1327,SI1328,SI1329,SI1330,SI1331,SI1332,SI1333,SI1334,SI1335,SI1336,SI1337,SI1338,SI1339,SI1340,SI1341,SI1342,SI1343,SI1344,SI1345,SI1346,SI1347,SI1348,SI1349,SI1350,SI1351,SI1352,SI1353,SI1354,SI1355,SI1356,SI1357,SI1358,SI1359,SI1360,SI1361,SI1362,SI1363,SI1364,SI1365,SI1366,SI1367,SI1368,SI1369,SI1370,SI1371,SI1372,SI1373,SI1374,SI1375,SI1376,SI1377,SI1378,SI1379,SI1380,SI1381,SI1382,SI1383,SI1384,SI1385,SI1386,SI1387,SI1388,SI1389,SI1390,SI1391,SI1392,SI1393,SI1394,SI1395,SI1396,SI1397,SI1398,SI1399,SI1400,SI1401,SI1402,SI1403,SI1404,SI1405,SI1406,SI1407,SI1408,SI1409,SI1410,SI1411,SI1412,SI1413,SI1414,SI1415,SI1416,SI1417,SI1418,SI1419,SI1420,SI1421,SI1422,SI1423,SI1424,SI1425,SI1426,SI1427,SI1428,SI1429,SI1430,SI1431,SI1432,SI1433,SI1434,SI1435,SI1436,SI1437,SI1438,SI1439,SI1440,SI1441,SI1442,SI1443,SI1444,SI1445,SI1446,SI1447,SI1448,SI1449,SI1450,SI1451,SI1452,SI1453,SI1454,SI1455,SI1456,SI1457,SI1458,SI1459,SI1460,SI1461,SI1462,SI1463,SI1464,SI1465,SI1466,SI1467,SI1468,SI1469,SI1470,SI1471,SI1472,SI1473,SI1474,SI1475,SI1476,SI1477,SI1478,SI1479,SI1480,SI1481,SI1482,SI1483,SI1484,SI1485,SI1486,SI1487,SI1488,SI1489,SI1490,SI1491,SI1492,SI1493,SI1494,SI1495,SI1496,SI1497,SI1498,SI1499,SI1500,SI1501,SI1502,SI1503,SI1504,SI1505,SI1506,SI1507,SI1508,SI1509,SI1510,SI1511,SI1512,SI1513,SI1514,SI1515,SI1516,SI1517,SI1518,SI1519,SI1520,SI1521,SI1522,SI1523,SI1524,SI1525,SI1526,SI1527,SI1528,SI1529,SI1530,SI1531,SI1532,SI1533,SI1534,SI1535,SI1536,SI1537,SI1538,SI1539,SI1540,SI1541,SI1542,SI1543,SI1544,SI1545,SI1546,SI1547,SI1548,SI1549,SI1550,SI1551,SI1552,SI1553,SI1554,SI1555,SI1556,SI1557,SI1558,SI1559,SI1560,SI1561,SI1562,SI1563,SI1564,SI1565,SI1566,SI1567,SI1568,SI1569,SI1570,SI1571,SI1572,SI1573,SI1574,SI1575,SI1576,SI1577,SI1578,SI1579,SI1580,SI1581,SI1582,SI1583,SI1584,SI1585,SI1586,SI1587,SI1588,SI1589,SI1590,SI1591,SI1592,SI1593,SI1594,SI1595,SI1596,SI1597,SI1598,SI1599,SI1600,SI1601,SI1602,SI1603,SI1604,SI1605,SI1606,SI1607,SI1608,SI1609,SI1610,SI1611,SI1612,SI1613,SI1614,SI1615,SI1616,SI1617,SI1618,SI1619,SI1620,SI1621,SI1622,SI1623,SI1624,SI1625,SI1626,SI1627,SI1628,SI1629,SI1630,SI1631,SI1632,SI1633,SI1634,SI1635,SI1636,SI1637,SI1638,SI1639,SI1640,SI1641,SI1642,SI1643,SI1644,SI1645,SI1646,SI1647,SI1648,SI1649,SI1650,SI1651,SI1652,SI1653,SI1654,SI1655,SI1656,SI1657,SI1658,SI1659,SI1660,SI1661,SI1662,SI1663,SI1664,SI1665,SI1666,SI1667,SI1668,SI1669,SI1670,SI1671,SI1672,SI1673,SI1674,SI1675,SI1676,SI1677,SI1678,SI1679,SI1680,SI1681,SI1682,SI1683,SI1684,SI1685,SI1686,SI1687,SI1688,SI1689,SI1690,SI1691,SI1692,SI1693,SI1694,SI1695,SI1696,SI1697,SI1698,SI1699,SI1700,SI1701,SI1702,SI1703,SI1704,SI1705,SI1706,SI1707,SI1708,SI1709,SI1710,SI1711,SI1712,SI1713,SI1714,SI1715,SI1716,SI1717,SI1718,SI1719,SI1720,SI1721,SI1722,SI1723,SI1724,SI1725,SI1726,SI1727,SI1728,SI1729,SI1730,SI1731,SI1732,SI1733,SI1734,SI1735,SI1736,SI1737,SI1738,SI1739,SI1740,SI1741,SI1742,SI1743,SI1744,SI1745,SI1746,SI1747,SI1748,SI1749,SI1750,SI1751,SI1752,SI1753,SI1754,SI1755,SI1756,SI1757,SI1758,SI1759,SI1760,SI1761,SI1762,SI1763,SI1764,SI1765,SI1766,SI1767,SI1768,SI1769,SI1770,SI1771,SI1772,SI1773,SI1774,SI1775,SI1776,SI1777,SI1778,SI1779,SI1780,SI1781,SI1782,SI1783,SI1784,SI1785,SI1786,SI1787,SI1788,SI1789,SI1790,SI1791,SI1792,SI1793,SI1794,SI1795,SI1796,SI1797,SI1798,SI1799,SI1800,SI1801,SI1802,SI1803,SI1804,SI1805,SI1806,SI1807,SI1808,SI1809,SI1810,SI1811,SI1812,SI1813,SI1814,SI1815,SI1816,SI1817,SI1818,SI1819,SI1820,SI1821,SI1822,SI1823,SI1824,SI1825,SI1826,SI1827,SI1828,SI1829,SI1830,SI1831,SI1832,SI1833,SI1834,SI1835,SI1836,SI1837,SI1838,SI1839,SI1840,SI1841,SI1842,SI1843,SI1844,SI1845,SI1846,SI1847,SI1848,SI1849,SI1850,SI1851,SI1852,SI1853,SI1854,SI1855,SI1856,SI1857,SI1858,SI1859,SI1860,SI1861,SI1862,SI1863,SI1864,SI1865,SI1866,SI1867,SI1868,SI1869,SI1870,SI1871,SI1872,SI1873,SI1874,SI1875,SI1876,SI1877,SI1878,SI1879,SI1880,SI1881,SI1882,SI1883,SI1884,SI1885,SI1886,SI1887,SI1888,SI1889,SI1890,SI1891,SI1892,SI1893,SI1894,SI1895,SI1896,SI1897,SI1898,SI1899,SI1900,SI1901,SI1902,SI1903,SI1904,SI1905,SI1906,SI1907,SI1908,SI1909,SI1910,SI1911,SI1912,SI1913,SI1914,SI1915,SI1916,SI1917,SI1918,SI1919,SI1920,SI1921,SI1922,SI1923,SI1924,SI1925,SI1926,SI1927,SI1928,SI1929,SI1930,SI1931,SI1932,SI1933,SI1934,SI1935,SI1936,SI1937,SI1938,SI1939,SI1940,SI1941,SI1942,SI1943,SI1944,SI1945,SI1946,SI1947,SI1948,SI1949,SI1950,SI1951,SI1952,SI1953,SI1954,SI1955,SI1956,SI1957,SI1958,SI1959,SI1960,SI1961,SI1962,SI1963,SI1964,SI1965,SI1966,SI1967,SI1968,SI1969,SI1970,SI1971,SI1972,SI1973,SI1974,SI1975,SI1976,SI1977,SI1978,SI1979,SI1980,SI1981,SI1982,SI1983,SI1984,SI1985,SI1986,SI1987,SI1988,SI1989,SI1990,SI1991,SI1992,SI1993,SI1994,SI1995,SI1996,SI1997,SI1998,SI1999,SI2000,SI2001,SI2002,SI2003,SI2004,SI2005,SI2006,SI2007,SI2008,SI2009,SI2010,SI2011,SI2012,SI2013,SI2014,SI2015,SI2016,SI2017,SI2018,SI2019,SI2020,SI2021,SI2022,SI2023,SI2024,SI2025,SI2026,SI2027,SI2028,SI2029,SI2030,SI2031,SI2032,SI2033,SI2034,SI2035,SI2036,SI2037,SI2038,SI2039,SI2040,SI2041,SI2042,SI2043,SI2044,SI2045,SI2046,SI2047,SI2048,SI2049,SI2050,SI2051,SI2052,SI2053,SI2054,SI2055,SI2056,SI2057,SI2058,SI2059,SI2060,SI2061,SI2062,SI2063,SI2064,SI2065,SI2066,SI2067,SI2068,SI2069,SI2070,SI2071,SI2072,SI2073,SI2074,SI2075,SI2076,SI2077,SI2078,SI2079,SI2080,SI2081,SI2082,SI2083,SI2084,SI2085,SI2086,SI2087,SI2088,SI2089,SI2090,SI2091,SI2092,SI2093,SI2094,SI2095,SI2096,SI2097,SI2098,SI2099,SI2100,SI2101,SI2102,SI2103,SI2104,SI2105,SI2106,SI2107,SI2108,SI2109,SI2110,SI2111,SI2112,SI2113,SI2114,SI2115,SI2116,SI2117,SI2118,SI2119,SI2120,SI2121,SI2122,SI2123,SI2124,SI2125,SI2126,SI2127,SI2128,SI2129,SI2130,SI2131,SI2132,SI2133,SI2134,SI2135,SI2136,SI2137,SI2138,SI2139,SI2140,SI2141,SI2142,SI2143,SI2144,SI2145,SI2146,SI2147,SI2148,SI2149,SI2150,SI2151,SI2152,SI2153,SI2154,SI2155,SI2156,SI2157,SI2158,SI2159,SI2160,SI2161,SI2162,SI2163,SI2164,SI2165,SI2166,SI2167,SI2168,SI2169,SI2170,SI2171,SI2172,SI2173,SI2174,SI2175,SI2176,SI2177,SI2178,SI2179,SI2180,SI2181,SI2182,SI2183,SI2184,SI2185,SI2186,SI2187,SI2188,SI2189,SI2190,SI2191,SI2192,SI2193,SI2194,SI2195,SI2196,SI2197,SI2198,SI2199,SI2200,SI2201,SI2202,SI2203,SI2204,SI2205,SI2206,SI2207,SI2208,SI2209,SI2210,SI2211,SI2212,SI2213,SI2214,SI2215,SI2216,SI2217,SI2218,SI2219,SI2220,SI2221,SI2222,SI2223,SI2224,SI2225,SI2226,SI2227,SI2228,SI2229,SI2230,SI2231,SI2232,SI2233,SI2234,SI2235,SI2236,SI2237,SI2238,SI2239,SI2240,SI2241,SI2242,SI2243,SI2244,SI2245,SI2246,SI2247,SI2248,SI2249,SI2250,SI2251,SI2252,SI2253,SI2254,SI2255,SI2256,SI2257,SI2258,SI2259,SI2260,SI2261,SI2262,SI2263,SI2264,SI2265,SI2266,SI2267,SI2268,SI2269,SI2270,SI2271,SI2272,SI2273,SI2274,SI2275,SI2276,SI2277,SI2278,SI2279,SI2280,SI2281,SI2282,SI2283,SI2284,SI2285,SI2286,SI2287,SI2288,SI2289,SI2290,SI2291,SI2292,SI2293,SI2294,SI2295,SI2296,SI2297,SI2298,SI2299,SI2300,SI2301,SI2302,SI2303,SI2304:std_logic;
signal end_vn1,end_vn2,end_vn3,end_vn4,end_vn5,end_vn6,end_vn7,end_vn8,end_vn9,end_vn10,end_vn11,end_vn12,end_vn13,end_vn14,end_vn15,end_vn16,end_vn17,end_vn18,end_vn19,end_vn20,end_vn21,end_vn22,end_vn23,end_vn24,end_vn25,end_vn26,end_vn27,end_vn28,end_vn29,end_vn30,end_vn31,end_vn32,end_vn33,end_vn34,end_vn35,end_vn36,end_vn37,end_vn38,end_vn39,end_vn40,end_vn41,end_vn42,end_vn43,end_vn44,end_vn45,end_vn46,end_vn47,end_vn48,end_vn49,end_vn50,end_vn51,end_vn52,end_vn53,end_vn54,end_vn55,end_vn56,end_vn57,end_vn58,end_vn59,end_vn60,end_vn61,end_vn62,end_vn63,end_vn64,end_vn65,end_vn66,end_vn67,end_vn68,end_vn69,end_vn70,end_vn71,end_vn72,end_vn73,end_vn74,end_vn75,end_vn76,end_vn77,end_vn78,end_vn79,end_vn80,end_vn81,end_vn82,end_vn83,end_vn84,end_vn85,end_vn86,end_vn87,end_vn88,end_vn89,end_vn90,end_vn91,end_vn92,end_vn93,end_vn94,end_vn95,end_vn96,end_vn97,end_vn98,end_vn99,end_vn100,end_vn101,end_vn102,end_vn103,end_vn104,end_vn105,end_vn106,end_vn107,end_vn108,end_vn109,end_vn110,end_vn111,end_vn112,end_vn113,end_vn114,end_vn115,end_vn116,end_vn117,end_vn118,end_vn119,end_vn120,end_vn121,end_vn122,end_vn123,end_vn124,end_vn125,end_vn126,end_vn127,end_vn128,end_vn129,end_vn130,end_vn131,end_vn132,end_vn133,end_vn134,end_vn135,end_vn136,end_vn137,end_vn138,end_vn139,end_vn140,end_vn141,end_vn142,end_vn143,end_vn144,end_vn145,end_vn146,end_vn147,end_vn148,end_vn149,end_vn150,end_vn151,end_vn152,end_vn153,end_vn154,end_vn155,end_vn156,end_vn157,end_vn158,end_vn159,end_vn160,end_vn161,end_vn162,end_vn163,end_vn164,end_vn165,end_vn166,end_vn167,end_vn168,end_vn169,end_vn170,end_vn171,end_vn172,end_vn173,end_vn174,end_vn175,end_vn176,end_vn177,end_vn178,end_vn179,end_vn180,end_vn181,end_vn182,end_vn183,end_vn184,end_vn185,end_vn186,end_vn187,end_vn188,end_vn189,end_vn190,end_vn191,end_vn192,end_vn193,end_vn194,end_vn195,end_vn196,end_vn197,end_vn198,end_vn199,end_vn200,end_vn201,end_vn202,end_vn203,end_vn204,end_vn205,end_vn206,end_vn207,end_vn208,end_vn209,end_vn210,end_vn211,end_vn212,end_vn213,end_vn214,end_vn215,end_vn216,end_vn217,end_vn218,end_vn219,end_vn220,end_vn221,end_vn222,end_vn223,end_vn224,end_vn225,end_vn226,end_vn227,end_vn228,end_vn229,end_vn230,end_vn231,end_vn232,end_vn233,end_vn234,end_vn235,end_vn236,end_vn237,end_vn238,end_vn239,end_vn240,end_vn241,end_vn242,end_vn243,end_vn244,end_vn245,end_vn246,end_vn247,end_vn248,end_vn249,end_vn250,end_vn251,end_vn252,end_vn253,end_vn254,end_vn255,end_vn256,end_vn257,end_vn258,end_vn259,end_vn260,end_vn261,end_vn262,end_vn263,end_vn264,end_vn265,end_vn266,end_vn267,end_vn268,end_vn269,end_vn270,end_vn271,end_vn272,end_vn273,end_vn274,end_vn275,end_vn276,end_vn277,end_vn278,end_vn279,end_vn280,end_vn281,end_vn282,end_vn283,end_vn284,end_vn285,end_vn286,end_vn287,end_vn288,end_vn289,end_vn290,end_vn291,end_vn292,end_vn293,end_vn294,end_vn295,end_vn296,end_vn297,end_vn298,end_vn299,end_vn300,end_vn301,end_vn302,end_vn303,end_vn304,end_vn305,end_vn306,end_vn307,end_vn308,end_vn309,end_vn310,end_vn311,end_vn312,end_vn313,end_vn314,end_vn315,end_vn316,end_vn317,end_vn318,end_vn319,end_vn320,end_vn321,end_vn322,end_vn323,end_vn324,end_vn325,end_vn326,end_vn327,end_vn328,end_vn329,end_vn330,end_vn331,end_vn332,end_vn333,end_vn334,end_vn335,end_vn336,end_vn337,end_vn338,end_vn339,end_vn340,end_vn341,end_vn342,end_vn343,end_vn344,end_vn345,end_vn346,end_vn347,end_vn348,end_vn349,end_vn350,end_vn351,end_vn352,end_vn353,end_vn354,end_vn355,end_vn356,end_vn357,end_vn358,end_vn359,end_vn360,end_vn361,end_vn362,end_vn363,end_vn364,end_vn365,end_vn366,end_vn367,end_vn368,end_vn369,end_vn370,end_vn371,end_vn372,end_vn373,end_vn374,end_vn375,end_vn376,end_vn377,end_vn378,end_vn379,end_vn380,end_vn381,end_vn382,end_vn383,end_vn384,end_vn385,end_vn386,end_vn387,end_vn388,end_vn389,end_vn390,end_vn391,end_vn392,end_vn393,end_vn394,end_vn395,end_vn396,end_vn397,end_vn398,end_vn399,end_vn400,end_vn401,end_vn402,end_vn403,end_vn404,end_vn405,end_vn406,end_vn407,end_vn408,end_vn409,end_vn410,end_vn411,end_vn412,end_vn413,end_vn414,end_vn415,end_vn416,end_vn417,end_vn418,end_vn419,end_vn420,end_vn421,end_vn422,end_vn423,end_vn424,end_vn425,end_vn426,end_vn427,end_vn428,end_vn429,end_vn430,end_vn431,end_vn432,end_vn433,end_vn434,end_vn435,end_vn436,end_vn437,end_vn438,end_vn439,end_vn440,end_vn441,end_vn442,end_vn443,end_vn444,end_vn445,end_vn446,end_vn447,end_vn448,end_vn449,end_vn450,end_vn451,end_vn452,end_vn453,end_vn454,end_vn455,end_vn456,end_vn457,end_vn458,end_vn459,end_vn460,end_vn461,end_vn462,end_vn463,end_vn464,end_vn465,end_vn466,end_vn467,end_vn468,end_vn469,end_vn470,end_vn471,end_vn472,end_vn473,end_vn474,end_vn475,end_vn476,end_vn477,end_vn478,end_vn479,end_vn480,end_vn481,end_vn482,end_vn483,end_vn484,end_vn485,end_vn486,end_vn487,end_vn488,end_vn489,end_vn490,end_vn491,end_vn492,end_vn493,end_vn494,end_vn495,end_vn496,end_vn497,end_vn498,end_vn499,end_vn500,end_vn501,end_vn502,end_vn503,end_vn504,end_vn505,end_vn506,end_vn507,end_vn508,end_vn509,end_vn510,end_vn511,end_vn512,end_vn513,end_vn514,end_vn515,end_vn516,end_vn517,end_vn518,end_vn519,end_vn520,end_vn521,end_vn522,end_vn523,end_vn524,end_vn525,end_vn526,end_vn527,end_vn528,end_vn529,end_vn530,end_vn531,end_vn532,end_vn533,end_vn534,end_vn535,end_vn536,end_vn537,end_vn538,end_vn539,end_vn540,end_vn541,end_vn542,end_vn543,end_vn544,end_vn545,end_vn546,end_vn547,end_vn548,end_vn549,end_vn550,end_vn551,end_vn552,end_vn553,end_vn554,end_vn555,end_vn556,end_vn557,end_vn558,end_vn559,end_vn560,end_vn561,end_vn562,end_vn563,end_vn564,end_vn565,end_vn566,end_vn567,end_vn568,end_vn569,end_vn570,end_vn571,end_vn572,end_vn573,end_vn574,end_vn575,end_vn576,end_vn577,end_vn578,end_vn579,end_vn580,end_vn581,end_vn582,end_vn583,end_vn584,end_vn585,end_vn586,end_vn587,end_vn588,end_vn589,end_vn590,end_vn591,end_vn592,end_vn593,end_vn594,end_vn595,end_vn596,end_vn597,end_vn598,end_vn599,end_vn600,end_vn601,end_vn602,end_vn603,end_vn604,end_vn605,end_vn606,end_vn607,end_vn608,end_vn609,end_vn610,end_vn611,end_vn612,end_vn613,end_vn614,end_vn615,end_vn616,end_vn617,end_vn618,end_vn619,end_vn620,end_vn621,end_vn622,end_vn623,end_vn624,end_vn625,end_vn626,end_vn627,end_vn628,end_vn629,end_vn630,end_vn631,end_vn632,end_vn633,end_vn634,end_vn635,end_vn636,end_vn637,end_vn638,end_vn639,end_vn640,end_vn641,end_vn642,end_vn643,end_vn644,end_vn645,end_vn646,end_vn647,end_vn648,end_vn649,end_vn650,end_vn651,end_vn652,end_vn653,end_vn654,end_vn655,end_vn656,end_vn657,end_vn658,end_vn659,end_vn660,end_vn661,end_vn662,end_vn663,end_vn664,end_vn665,end_vn666,end_vn667,end_vn668,end_vn669,end_vn670,end_vn671,end_vn672,end_vn673,end_vn674,end_vn675,end_vn676,end_vn677,end_vn678,end_vn679,end_vn680,end_vn681,end_vn682,end_vn683,end_vn684,end_vn685,end_vn686,end_vn687,end_vn688,end_vn689,end_vn690,end_vn691,end_vn692,end_vn693,end_vn694,end_vn695,end_vn696,end_vn697,end_vn698,end_vn699,end_vn700,end_vn701,end_vn702,end_vn703,end_vn704,end_vn705,end_vn706,end_vn707,end_vn708,end_vn709,end_vn710,end_vn711,end_vn712,end_vn713,end_vn714,end_vn715,end_vn716,end_vn717,end_vn718,end_vn719,end_vn720,end_vn721,end_vn722,end_vn723,end_vn724,end_vn725,end_vn726,end_vn727,end_vn728,end_vn729,end_vn730,end_vn731,end_vn732,end_vn733,end_vn734,end_vn735,end_vn736,end_vn737,end_vn738,end_vn739,end_vn740,end_vn741,end_vn742,end_vn743,end_vn744,end_vn745,end_vn746,end_vn747,end_vn748,end_vn749,end_vn750,end_vn751,end_vn752,end_vn753,end_vn754,end_vn755,end_vn756,end_vn757,end_vn758,end_vn759,end_vn760,end_vn761,end_vn762,end_vn763,end_vn764,end_vn765,end_vn766,end_vn767,end_vn768,end_vn769,end_vn770,end_vn771,end_vn772,end_vn773,end_vn774,end_vn775,end_vn776,end_vn777,end_vn778,end_vn779,end_vn780,end_vn781,end_vn782,end_vn783,end_vn784,end_vn785,end_vn786,end_vn787,end_vn788,end_vn789,end_vn790,end_vn791,end_vn792,end_vn793,end_vn794,end_vn795,end_vn796,end_vn797,end_vn798,end_vn799,end_vn800,end_vn801,end_vn802,end_vn803,end_vn804,end_vn805,end_vn806,end_vn807,end_vn808,end_vn809,end_vn810,end_vn811,end_vn812,end_vn813,end_vn814,end_vn815,end_vn816,end_vn817,end_vn818,end_vn819,end_vn820,end_vn821,end_vn822,end_vn823,end_vn824,end_vn825,end_vn826,end_vn827,end_vn828,end_vn829,end_vn830,end_vn831,end_vn832,end_vn833,end_vn834,end_vn835,end_vn836,end_vn837,end_vn838,end_vn839,end_vn840,end_vn841,end_vn842,end_vn843,end_vn844,end_vn845,end_vn846,end_vn847,end_vn848,end_vn849,end_vn850,end_vn851,end_vn852,end_vn853,end_vn854,end_vn855,end_vn856,end_vn857,end_vn858,end_vn859,end_vn860,end_vn861,end_vn862,end_vn863,end_vn864,end_vn865,end_vn866,end_vn867,end_vn868,end_vn869,end_vn870,end_vn871,end_vn872,end_vn873,end_vn874,end_vn875,end_vn876,end_vn877,end_vn878,end_vn879,end_vn880,end_vn881,end_vn882,end_vn883,end_vn884,end_vn885,end_vn886,end_vn887,end_vn888,end_vn889,end_vn890,end_vn891,end_vn892,end_vn893,end_vn894,end_vn895,end_vn896,end_vn897,end_vn898,end_vn899,end_vn900,end_vn901,end_vn902,end_vn903,end_vn904,end_vn905,end_vn906,end_vn907,end_vn908,end_vn909,end_vn910,end_vn911,end_vn912,end_vn913,end_vn914,end_vn915,end_vn916,end_vn917,end_vn918,end_vn919,end_vn920,end_vn921,end_vn922,end_vn923,end_vn924,end_vn925,end_vn926,end_vn927,end_vn928,end_vn929,end_vn930,end_vn931,end_vn932,end_vn933,end_vn934,end_vn935,end_vn936,end_vn937,end_vn938,end_vn939,end_vn940,end_vn941,end_vn942,end_vn943,end_vn944,end_vn945,end_vn946,end_vn947,end_vn948,end_vn949,end_vn950,end_vn951,end_vn952,end_vn953,end_vn954,end_vn955,end_vn956,end_vn957,end_vn958,end_vn959,end_vn960,end_vn961,end_vn962,end_vn963,end_vn964,end_vn965,end_vn966,end_vn967,end_vn968,end_vn969,end_vn970,end_vn971,end_vn972,end_vn973,end_vn974,end_vn975,end_vn976,end_vn977,end_vn978,end_vn979,end_vn980,end_vn981,end_vn982,end_vn983,end_vn984,end_vn985,end_vn986,end_vn987,end_vn988,end_vn989,end_vn990,end_vn991,end_vn992,end_vn993,end_vn994,end_vn995,end_vn996,end_vn997,end_vn998,end_vn999,end_vn1000,end_vn1001,end_vn1002,end_vn1003,end_vn1004,end_vn1005,end_vn1006,end_vn1007,end_vn1008,end_vn1009,end_vn1010,end_vn1011,end_vn1012,end_vn1013,end_vn1014,end_vn1015,end_vn1016,end_vn1017,end_vn1018,end_vn1019,end_vn1020,end_vn1021,end_vn1022,end_vn1023,end_vn1024,end_vn1025,end_vn1026,end_vn1027,end_vn1028,end_vn1029,end_vn1030,end_vn1031,end_vn1032,end_vn1033,end_vn1034,end_vn1035,end_vn1036,end_vn1037,end_vn1038,end_vn1039,end_vn1040,end_vn1041,end_vn1042,end_vn1043,end_vn1044,end_vn1045,end_vn1046,end_vn1047,end_vn1048,end_vn1049,end_vn1050,end_vn1051,end_vn1052,end_vn1053,end_vn1054,end_vn1055,end_vn1056,end_vn1057,end_vn1058,end_vn1059,end_vn1060,end_vn1061,end_vn1062,end_vn1063,end_vn1064,end_vn1065,end_vn1066,end_vn1067,end_vn1068,end_vn1069,end_vn1070,end_vn1071,end_vn1072,end_vn1073,end_vn1074,end_vn1075,end_vn1076,end_vn1077,end_vn1078,end_vn1079,end_vn1080,end_vn1081,end_vn1082,end_vn1083,end_vn1084,end_vn1085,end_vn1086,end_vn1087,end_vn1088,end_vn1089,end_vn1090,end_vn1091,end_vn1092,end_vn1093,end_vn1094,end_vn1095,end_vn1096,end_vn1097,end_vn1098,end_vn1099,end_vn1100,end_vn1101,end_vn1102,end_vn1103,end_vn1104,end_vn1105,end_vn1106,end_vn1107,end_vn1108,end_vn1109,end_vn1110,end_vn1111,end_vn1112,end_vn1113,end_vn1114,end_vn1115,end_vn1116,end_vn1117,end_vn1118,end_vn1119,end_vn1120,end_vn1121,end_vn1122,end_vn1123,end_vn1124,end_vn1125,end_vn1126,end_vn1127,end_vn1128,end_vn1129,end_vn1130,end_vn1131,end_vn1132,end_vn1133,end_vn1134,end_vn1135,end_vn1136,end_vn1137,end_vn1138,end_vn1139,end_vn1140,end_vn1141,end_vn1142,end_vn1143,end_vn1144,end_vn1145,end_vn1146,end_vn1147,end_vn1148,end_vn1149,end_vn1150,end_vn1151,end_vn1152,end_vn1153,end_vn1154,end_vn1155,end_vn1156,end_vn1157,end_vn1158,end_vn1159,end_vn1160,end_vn1161,end_vn1162,end_vn1163,end_vn1164,end_vn1165,end_vn1166,end_vn1167,end_vn1168,end_vn1169,end_vn1170,end_vn1171,end_vn1172,end_vn1173,end_vn1174,end_vn1175,end_vn1176,end_vn1177,end_vn1178,end_vn1179,end_vn1180,end_vn1181,end_vn1182,end_vn1183,end_vn1184,end_vn1185,end_vn1186,end_vn1187,end_vn1188,end_vn1189,end_vn1190,end_vn1191,end_vn1192,end_vn1193,end_vn1194,end_vn1195,end_vn1196,end_vn1197,end_vn1198,end_vn1199,end_vn1200,end_vn1201,end_vn1202,end_vn1203,end_vn1204,end_vn1205,end_vn1206,end_vn1207,end_vn1208,end_vn1209,end_vn1210,end_vn1211,end_vn1212,end_vn1213,end_vn1214,end_vn1215,end_vn1216,end_vn1217,end_vn1218,end_vn1219,end_vn1220,end_vn1221,end_vn1222,end_vn1223,end_vn1224,end_vn1225,end_vn1226,end_vn1227,end_vn1228,end_vn1229,end_vn1230,end_vn1231,end_vn1232,end_vn1233,end_vn1234,end_vn1235,end_vn1236,end_vn1237,end_vn1238,end_vn1239,end_vn1240,end_vn1241,end_vn1242,end_vn1243,end_vn1244,end_vn1245,end_vn1246,end_vn1247,end_vn1248,end_vn1249,end_vn1250,end_vn1251,end_vn1252,end_vn1253,end_vn1254,end_vn1255,end_vn1256,end_vn1257,end_vn1258,end_vn1259,end_vn1260,end_vn1261,end_vn1262,end_vn1263,end_vn1264,end_vn1265,end_vn1266,end_vn1267,end_vn1268,end_vn1269,end_vn1270,end_vn1271,end_vn1272,end_vn1273,end_vn1274,end_vn1275,end_vn1276,end_vn1277,end_vn1278,end_vn1279,end_vn1280,end_vn1281,end_vn1282,end_vn1283,end_vn1284,end_vn1285,end_vn1286,end_vn1287,end_vn1288,end_vn1289,end_vn1290,end_vn1291,end_vn1292,end_vn1293,end_vn1294,end_vn1295,end_vn1296,end_vn1297,end_vn1298,end_vn1299,end_vn1300,end_vn1301,end_vn1302,end_vn1303,end_vn1304,end_vn1305,end_vn1306,end_vn1307,end_vn1308,end_vn1309,end_vn1310,end_vn1311,end_vn1312,end_vn1313,end_vn1314,end_vn1315,end_vn1316,end_vn1317,end_vn1318,end_vn1319,end_vn1320,end_vn1321,end_vn1322,end_vn1323,end_vn1324,end_vn1325,end_vn1326,end_vn1327,end_vn1328,end_vn1329,end_vn1330,end_vn1331,end_vn1332,end_vn1333,end_vn1334,end_vn1335,end_vn1336,end_vn1337,end_vn1338,end_vn1339,end_vn1340,end_vn1341,end_vn1342,end_vn1343,end_vn1344,end_vn1345,end_vn1346,end_vn1347,end_vn1348,end_vn1349,end_vn1350,end_vn1351,end_vn1352,end_vn1353,end_vn1354,end_vn1355,end_vn1356,end_vn1357,end_vn1358,end_vn1359,end_vn1360,end_vn1361,end_vn1362,end_vn1363,end_vn1364,end_vn1365,end_vn1366,end_vn1367,end_vn1368,end_vn1369,end_vn1370,end_vn1371,end_vn1372,end_vn1373,end_vn1374,end_vn1375,end_vn1376,end_vn1377,end_vn1378,end_vn1379,end_vn1380,end_vn1381,end_vn1382,end_vn1383,end_vn1384,end_vn1385,end_vn1386,end_vn1387,end_vn1388,end_vn1389,end_vn1390,end_vn1391,end_vn1392,end_vn1393,end_vn1394,end_vn1395,end_vn1396,end_vn1397,end_vn1398,end_vn1399,end_vn1400,end_vn1401,end_vn1402,end_vn1403,end_vn1404,end_vn1405,end_vn1406,end_vn1407,end_vn1408,end_vn1409,end_vn1410,end_vn1411,end_vn1412,end_vn1413,end_vn1414,end_vn1415,end_vn1416,end_vn1417,end_vn1418,end_vn1419,end_vn1420,end_vn1421,end_vn1422,end_vn1423,end_vn1424,end_vn1425,end_vn1426,end_vn1427,end_vn1428,end_vn1429,end_vn1430,end_vn1431,end_vn1432,end_vn1433,end_vn1434,end_vn1435,end_vn1436,end_vn1437,end_vn1438,end_vn1439,end_vn1440,end_vn1441,end_vn1442,end_vn1443,end_vn1444,end_vn1445,end_vn1446,end_vn1447,end_vn1448,end_vn1449,end_vn1450,end_vn1451,end_vn1452,end_vn1453,end_vn1454,end_vn1455,end_vn1456,end_vn1457,end_vn1458,end_vn1459,end_vn1460,end_vn1461,end_vn1462,end_vn1463,end_vn1464,end_vn1465,end_vn1466,end_vn1467,end_vn1468,end_vn1469,end_vn1470,end_vn1471,end_vn1472,end_vn1473,end_vn1474,end_vn1475,end_vn1476,end_vn1477,end_vn1478,end_vn1479,end_vn1480,end_vn1481,end_vn1482,end_vn1483,end_vn1484,end_vn1485,end_vn1486,end_vn1487,end_vn1488,end_vn1489,end_vn1490,end_vn1491,end_vn1492,end_vn1493,end_vn1494,end_vn1495,end_vn1496,end_vn1497,end_vn1498,end_vn1499,end_vn1500,end_vn1501,end_vn1502,end_vn1503,end_vn1504,end_vn1505,end_vn1506,end_vn1507,end_vn1508,end_vn1509,end_vn1510,end_vn1511,end_vn1512,end_vn1513,end_vn1514,end_vn1515,end_vn1516,end_vn1517,end_vn1518,end_vn1519,end_vn1520,end_vn1521,end_vn1522,end_vn1523,end_vn1524,end_vn1525,end_vn1526,end_vn1527,end_vn1528,end_vn1529,end_vn1530,end_vn1531,end_vn1532,end_vn1533,end_vn1534,end_vn1535,end_vn1536,end_vn1537,end_vn1538,end_vn1539,end_vn1540,end_vn1541,end_vn1542,end_vn1543,end_vn1544,end_vn1545,end_vn1546,end_vn1547,end_vn1548,end_vn1549,end_vn1550,end_vn1551,end_vn1552,end_vn1553,end_vn1554,end_vn1555,end_vn1556,end_vn1557,end_vn1558,end_vn1559,end_vn1560,end_vn1561,end_vn1562,end_vn1563,end_vn1564,end_vn1565,end_vn1566,end_vn1567,end_vn1568,end_vn1569,end_vn1570,end_vn1571,end_vn1572,end_vn1573,end_vn1574,end_vn1575,end_vn1576,end_vn1577,end_vn1578,end_vn1579,end_vn1580,end_vn1581,end_vn1582,end_vn1583,end_vn1584,end_vn1585,end_vn1586,end_vn1587,end_vn1588,end_vn1589,end_vn1590,end_vn1591,end_vn1592,end_vn1593,end_vn1594,end_vn1595,end_vn1596,end_vn1597,end_vn1598,end_vn1599,end_vn1600,end_vn1601,end_vn1602,end_vn1603,end_vn1604,end_vn1605,end_vn1606,end_vn1607,end_vn1608,end_vn1609,end_vn1610,end_vn1611,end_vn1612,end_vn1613,end_vn1614,end_vn1615,end_vn1616,end_vn1617,end_vn1618,end_vn1619,end_vn1620,end_vn1621,end_vn1622,end_vn1623,end_vn1624,end_vn1625,end_vn1626,end_vn1627,end_vn1628,end_vn1629,end_vn1630,end_vn1631,end_vn1632,end_vn1633,end_vn1634,end_vn1635,end_vn1636,end_vn1637,end_vn1638,end_vn1639,end_vn1640,end_vn1641,end_vn1642,end_vn1643,end_vn1644,end_vn1645,end_vn1646,end_vn1647,end_vn1648,end_vn1649,end_vn1650,end_vn1651,end_vn1652,end_vn1653,end_vn1654,end_vn1655,end_vn1656,end_vn1657,end_vn1658,end_vn1659,end_vn1660,end_vn1661,end_vn1662,end_vn1663,end_vn1664,end_vn1665,end_vn1666,end_vn1667,end_vn1668,end_vn1669,end_vn1670,end_vn1671,end_vn1672,end_vn1673,end_vn1674,end_vn1675,end_vn1676,end_vn1677,end_vn1678,end_vn1679,end_vn1680,end_vn1681,end_vn1682,end_vn1683,end_vn1684,end_vn1685,end_vn1686,end_vn1687,end_vn1688,end_vn1689,end_vn1690,end_vn1691,end_vn1692,end_vn1693,end_vn1694,end_vn1695,end_vn1696,end_vn1697,end_vn1698,end_vn1699,end_vn1700,end_vn1701,end_vn1702,end_vn1703,end_vn1704,end_vn1705,end_vn1706,end_vn1707,end_vn1708,end_vn1709,end_vn1710,end_vn1711,end_vn1712,end_vn1713,end_vn1714,end_vn1715,end_vn1716,end_vn1717,end_vn1718,end_vn1719,end_vn1720,end_vn1721,end_vn1722,end_vn1723,end_vn1724,end_vn1725,end_vn1726,end_vn1727,end_vn1728,end_vn1729,end_vn1730,end_vn1731,end_vn1732,end_vn1733,end_vn1734,end_vn1735,end_vn1736,end_vn1737,end_vn1738,end_vn1739,end_vn1740,end_vn1741,end_vn1742,end_vn1743,end_vn1744,end_vn1745,end_vn1746,end_vn1747,end_vn1748,end_vn1749,end_vn1750,end_vn1751,end_vn1752,end_vn1753,end_vn1754,end_vn1755,end_vn1756,end_vn1757,end_vn1758,end_vn1759,end_vn1760,end_vn1761,end_vn1762,end_vn1763,end_vn1764,end_vn1765,end_vn1766,end_vn1767,end_vn1768,end_vn1769,end_vn1770,end_vn1771,end_vn1772,end_vn1773,end_vn1774,end_vn1775,end_vn1776,end_vn1777,end_vn1778,end_vn1779,end_vn1780,end_vn1781,end_vn1782,end_vn1783,end_vn1784,end_vn1785,end_vn1786,end_vn1787,end_vn1788,end_vn1789,end_vn1790,end_vn1791,end_vn1792,end_vn1793,end_vn1794,end_vn1795,end_vn1796,end_vn1797,end_vn1798,end_vn1799,end_vn1800,end_vn1801,end_vn1802,end_vn1803,end_vn1804,end_vn1805,end_vn1806,end_vn1807,end_vn1808,end_vn1809,end_vn1810,end_vn1811,end_vn1812,end_vn1813,end_vn1814,end_vn1815,end_vn1816,end_vn1817,end_vn1818,end_vn1819,end_vn1820,end_vn1821,end_vn1822,end_vn1823,end_vn1824,end_vn1825,end_vn1826,end_vn1827,end_vn1828,end_vn1829,end_vn1830,end_vn1831,end_vn1832,end_vn1833,end_vn1834,end_vn1835,end_vn1836,end_vn1837,end_vn1838,end_vn1839,end_vn1840,end_vn1841,end_vn1842,end_vn1843,end_vn1844,end_vn1845,end_vn1846,end_vn1847,end_vn1848,end_vn1849,end_vn1850,end_vn1851,end_vn1852,end_vn1853,end_vn1854,end_vn1855,end_vn1856,end_vn1857,end_vn1858,end_vn1859,end_vn1860,end_vn1861,end_vn1862,end_vn1863,end_vn1864,end_vn1865,end_vn1866,end_vn1867,end_vn1868,end_vn1869,end_vn1870,end_vn1871,end_vn1872,end_vn1873,end_vn1874,end_vn1875,end_vn1876,end_vn1877,end_vn1878,end_vn1879,end_vn1880,end_vn1881,end_vn1882,end_vn1883,end_vn1884,end_vn1885,end_vn1886,end_vn1887,end_vn1888,end_vn1889,end_vn1890,end_vn1891,end_vn1892,end_vn1893,end_vn1894,end_vn1895,end_vn1896,end_vn1897,end_vn1898,end_vn1899,end_vn1900,end_vn1901,end_vn1902,end_vn1903,end_vn1904,end_vn1905,end_vn1906,end_vn1907,end_vn1908,end_vn1909,end_vn1910,end_vn1911,end_vn1912,end_vn1913,end_vn1914,end_vn1915,end_vn1916,end_vn1917,end_vn1918,end_vn1919,end_vn1920,end_vn1921,end_vn1922,end_vn1923,end_vn1924,end_vn1925,end_vn1926,end_vn1927,end_vn1928,end_vn1929,end_vn1930,end_vn1931,end_vn1932,end_vn1933,end_vn1934,end_vn1935,end_vn1936,end_vn1937,end_vn1938,end_vn1939,end_vn1940,end_vn1941,end_vn1942,end_vn1943,end_vn1944,end_vn1945,end_vn1946,end_vn1947,end_vn1948,end_vn1949,end_vn1950,end_vn1951,end_vn1952,end_vn1953,end_vn1954,end_vn1955,end_vn1956,end_vn1957,end_vn1958,end_vn1959,end_vn1960,end_vn1961,end_vn1962,end_vn1963,end_vn1964,end_vn1965,end_vn1966,end_vn1967,end_vn1968,end_vn1969,end_vn1970,end_vn1971,end_vn1972,end_vn1973,end_vn1974,end_vn1975,end_vn1976,end_vn1977,end_vn1978,end_vn1979,end_vn1980,end_vn1981,end_vn1982,end_vn1983,end_vn1984,end_vn1985,end_vn1986,end_vn1987,end_vn1988,end_vn1989,end_vn1990,end_vn1991,end_vn1992,end_vn1993,end_vn1994,end_vn1995,end_vn1996,end_vn1997,end_vn1998,end_vn1999,end_vn2000,end_vn2001,end_vn2002,end_vn2003,end_vn2004,end_vn2005,end_vn2006,end_vn2007,end_vn2008,end_vn2009,end_vn2010,end_vn2011,end_vn2012,end_vn2013,end_vn2014,end_vn2015,end_vn2016,end_vn2017,end_vn2018,end_vn2019,end_vn2020,end_vn2021,end_vn2022,end_vn2023,end_vn2024,end_vn2025,end_vn2026,end_vn2027,end_vn2028,end_vn2029,end_vn2030,end_vn2031,end_vn2032,end_vn2033,end_vn2034,end_vn2035,end_vn2036,end_vn2037,end_vn2038,end_vn2039,end_vn2040,end_vn2041,end_vn2042,end_vn2043,end_vn2044,end_vn2045,end_vn2046,end_vn2047,end_vn2048,end_vn2049,end_vn2050,end_vn2051,end_vn2052,end_vn2053,end_vn2054,end_vn2055,end_vn2056,end_vn2057,end_vn2058,end_vn2059,end_vn2060,end_vn2061,end_vn2062,end_vn2063,end_vn2064,end_vn2065,end_vn2066,end_vn2067,end_vn2068,end_vn2069,end_vn2070,end_vn2071,end_vn2072,end_vn2073,end_vn2074,end_vn2075,end_vn2076,end_vn2077,end_vn2078,end_vn2079,end_vn2080,end_vn2081,end_vn2082,end_vn2083,end_vn2084,end_vn2085,end_vn2086,end_vn2087,end_vn2088,end_vn2089,end_vn2090,end_vn2091,end_vn2092,end_vn2093,end_vn2094,end_vn2095,end_vn2096,end_vn2097,end_vn2098,end_vn2099,end_vn2100,end_vn2101,end_vn2102,end_vn2103,end_vn2104,end_vn2105,end_vn2106,end_vn2107,end_vn2108,end_vn2109,end_vn2110,end_vn2111,end_vn2112,end_vn2113,end_vn2114,end_vn2115,end_vn2116,end_vn2117,end_vn2118,end_vn2119,end_vn2120,end_vn2121,end_vn2122,end_vn2123,end_vn2124,end_vn2125,end_vn2126,end_vn2127,end_vn2128,end_vn2129,end_vn2130,end_vn2131,end_vn2132,end_vn2133,end_vn2134,end_vn2135,end_vn2136,end_vn2137,end_vn2138,end_vn2139,end_vn2140,end_vn2141,end_vn2142,end_vn2143,end_vn2144,end_vn2145,end_vn2146,end_vn2147,end_vn2148,end_vn2149,end_vn2150,end_vn2151,end_vn2152,end_vn2153,end_vn2154,end_vn2155,end_vn2156,end_vn2157,end_vn2158,end_vn2159,end_vn2160,end_vn2161,end_vn2162,end_vn2163,end_vn2164,end_vn2165,end_vn2166,end_vn2167,end_vn2168,end_vn2169,end_vn2170,end_vn2171,end_vn2172,end_vn2173,end_vn2174,end_vn2175,end_vn2176,end_vn2177,end_vn2178,end_vn2179,end_vn2180,end_vn2181,end_vn2182,end_vn2183,end_vn2184,end_vn2185,end_vn2186,end_vn2187,end_vn2188,end_vn2189,end_vn2190,end_vn2191,end_vn2192,end_vn2193,end_vn2194,end_vn2195,end_vn2196,end_vn2197,end_vn2198,end_vn2199,end_vn2200,end_vn2201,end_vn2202,end_vn2203,end_vn2204,end_vn2205,end_vn2206,end_vn2207,end_vn2208,end_vn2209,end_vn2210,end_vn2211,end_vn2212,end_vn2213,end_vn2214,end_vn2215,end_vn2216,end_vn2217,end_vn2218,end_vn2219,end_vn2220,end_vn2221,end_vn2222,end_vn2223,end_vn2224,end_vn2225,end_vn2226,end_vn2227,end_vn2228,end_vn2229,end_vn2230,end_vn2231,end_vn2232,end_vn2233,end_vn2234,end_vn2235,end_vn2236,end_vn2237,end_vn2238,end_vn2239,end_vn2240,end_vn2241,end_vn2242,end_vn2243,end_vn2244,end_vn2245,end_vn2246,end_vn2247,end_vn2248,end_vn2249,end_vn2250,end_vn2251,end_vn2252,end_vn2253,end_vn2254,end_vn2255,end_vn2256,end_vn2257,end_vn2258,end_vn2259,end_vn2260,end_vn2261,end_vn2262,end_vn2263,end_vn2264,end_vn2265,end_vn2266,end_vn2267,end_vn2268,end_vn2269,end_vn2270,end_vn2271,end_vn2272,end_vn2273,end_vn2274,end_vn2275,end_vn2276,end_vn2277,end_vn2278,end_vn2279,end_vn2280,end_vn2281,end_vn2282,end_vn2283,end_vn2284,end_vn2285,end_vn2286,end_vn2287,end_vn2288,end_vn2289,end_vn2290,end_vn2291,end_vn2292,end_vn2293,end_vn2294,end_vn2295,end_vn2296,end_vn2297,end_vn2298,end_vn2299,end_vn2300,end_vn2301,end_vn2302,end_vn2303,end_vn2304:std_logic;
signal end_cn1,end_cn2,end_cn3,end_cn4,end_cn5,end_cn6,end_cn7,end_cn8,end_cn9,end_cn10,end_cn11,end_cn12,end_cn13,end_cn14,end_cn15,end_cn16,end_cn17,end_cn18,end_cn19,end_cn20,end_cn21,end_cn22,end_cn23,end_cn24,end_cn25,end_cn26,end_cn27,end_cn28,end_cn29,end_cn30,end_cn31,end_cn32,end_cn33,end_cn34,end_cn35,end_cn36,end_cn37,end_cn38,end_cn39,end_cn40,end_cn41,end_cn42,end_cn43,end_cn44,end_cn45,end_cn46,end_cn47,end_cn48,end_cn49,end_cn50,end_cn51,end_cn52,end_cn53,end_cn54,end_cn55,end_cn56,end_cn57,end_cn58,end_cn59,end_cn60,end_cn61,end_cn62,end_cn63,end_cn64,end_cn65,end_cn66,end_cn67,end_cn68,end_cn69,end_cn70,end_cn71,end_cn72,end_cn73,end_cn74,end_cn75,end_cn76,end_cn77,end_cn78,end_cn79,end_cn80,end_cn81,end_cn82,end_cn83,end_cn84,end_cn85,end_cn86,end_cn87,end_cn88,end_cn89,end_cn90,end_cn91,end_cn92,end_cn93,end_cn94,end_cn95,end_cn96,end_cn97,end_cn98,end_cn99,end_cn100,end_cn101,end_cn102,end_cn103,end_cn104,end_cn105,end_cn106,end_cn107,end_cn108,end_cn109,end_cn110,end_cn111,end_cn112,end_cn113,end_cn114,end_cn115,end_cn116,end_cn117,end_cn118,end_cn119,end_cn120,end_cn121,end_cn122,end_cn123,end_cn124,end_cn125,end_cn126,end_cn127,end_cn128,end_cn129,end_cn130,end_cn131,end_cn132,end_cn133,end_cn134,end_cn135,end_cn136,end_cn137,end_cn138,end_cn139,end_cn140,end_cn141,end_cn142,end_cn143,end_cn144,end_cn145,end_cn146,end_cn147,end_cn148,end_cn149,end_cn150,end_cn151,end_cn152,end_cn153,end_cn154,end_cn155,end_cn156,end_cn157,end_cn158,end_cn159,end_cn160,end_cn161,end_cn162,end_cn163,end_cn164,end_cn165,end_cn166,end_cn167,end_cn168,end_cn169,end_cn170,end_cn171,end_cn172,end_cn173,end_cn174,end_cn175,end_cn176,end_cn177,end_cn178,end_cn179,end_cn180,end_cn181,end_cn182,end_cn183,end_cn184,end_cn185,end_cn186,end_cn187,end_cn188,end_cn189,end_cn190,end_cn191,end_cn192,end_cn193,end_cn194,end_cn195,end_cn196,end_cn197,end_cn198,end_cn199,end_cn200,end_cn201,end_cn202,end_cn203,end_cn204,end_cn205,end_cn206,end_cn207,end_cn208,end_cn209,end_cn210,end_cn211,end_cn212,end_cn213,end_cn214,end_cn215,end_cn216,end_cn217,end_cn218,end_cn219,end_cn220,end_cn221,end_cn222,end_cn223,end_cn224,end_cn225,end_cn226,end_cn227,end_cn228,end_cn229,end_cn230,end_cn231,end_cn232,end_cn233,end_cn234,end_cn235,end_cn236,end_cn237,end_cn238,end_cn239,end_cn240,end_cn241,end_cn242,end_cn243,end_cn244,end_cn245,end_cn246,end_cn247,end_cn248,end_cn249,end_cn250,end_cn251,end_cn252,end_cn253,end_cn254,end_cn255,end_cn256,end_cn257,end_cn258,end_cn259,end_cn260,end_cn261,end_cn262,end_cn263,end_cn264,end_cn265,end_cn266,end_cn267,end_cn268,end_cn269,end_cn270,end_cn271,end_cn272,end_cn273,end_cn274,end_cn275,end_cn276,end_cn277,end_cn278,end_cn279,end_cn280,end_cn281,end_cn282,end_cn283,end_cn284,end_cn285,end_cn286,end_cn287,end_cn288,end_cn289,end_cn290,end_cn291,end_cn292,end_cn293,end_cn294,end_cn295,end_cn296,end_cn297,end_cn298,end_cn299,end_cn300,end_cn301,end_cn302,end_cn303,end_cn304,end_cn305,end_cn306,end_cn307,end_cn308,end_cn309,end_cn310,end_cn311,end_cn312,end_cn313,end_cn314,end_cn315,end_cn316,end_cn317,end_cn318,end_cn319,end_cn320,end_cn321,end_cn322,end_cn323,end_cn324,end_cn325,end_cn326,end_cn327,end_cn328,end_cn329,end_cn330,end_cn331,end_cn332,end_cn333,end_cn334,end_cn335,end_cn336,end_cn337,end_cn338,end_cn339,end_cn340,end_cn341,end_cn342,end_cn343,end_cn344,end_cn345,end_cn346,end_cn347,end_cn348,end_cn349,end_cn350,end_cn351,end_cn352,end_cn353,end_cn354,end_cn355,end_cn356,end_cn357,end_cn358,end_cn359,end_cn360,end_cn361,end_cn362,end_cn363,end_cn364,end_cn365,end_cn366,end_cn367,end_cn368,end_cn369,end_cn370,end_cn371,end_cn372,end_cn373,end_cn374,end_cn375,end_cn376,end_cn377,end_cn378,end_cn379,end_cn380,end_cn381,end_cn382,end_cn383,end_cn384,end_cn385,end_cn386,end_cn387,end_cn388,end_cn389,end_cn390,end_cn391,end_cn392,end_cn393,end_cn394,end_cn395,end_cn396,end_cn397,end_cn398,end_cn399,end_cn400,end_cn401,end_cn402,end_cn403,end_cn404,end_cn405,end_cn406,end_cn407,end_cn408,end_cn409,end_cn410,end_cn411,end_cn412,end_cn413,end_cn414,end_cn415,end_cn416,end_cn417,end_cn418,end_cn419,end_cn420,end_cn421,end_cn422,end_cn423,end_cn424,end_cn425,end_cn426,end_cn427,end_cn428,end_cn429,end_cn430,end_cn431,end_cn432,end_cn433,end_cn434,end_cn435,end_cn436,end_cn437,end_cn438,end_cn439,end_cn440,end_cn441,end_cn442,end_cn443,end_cn444,end_cn445,end_cn446,end_cn447,end_cn448,end_cn449,end_cn450,end_cn451,end_cn452,end_cn453,end_cn454,end_cn455,end_cn456,end_cn457,end_cn458,end_cn459,end_cn460,end_cn461,end_cn462,end_cn463,end_cn464,end_cn465,end_cn466,end_cn467,end_cn468,end_cn469,end_cn470,end_cn471,end_cn472,end_cn473,end_cn474,end_cn475,end_cn476,end_cn477,end_cn478,end_cn479,end_cn480,end_cn481,end_cn482,end_cn483,end_cn484,end_cn485,end_cn486,end_cn487,end_cn488,end_cn489,end_cn490,end_cn491,end_cn492,end_cn493,end_cn494,end_cn495,end_cn496,end_cn497,end_cn498,end_cn499,end_cn500,end_cn501,end_cn502,end_cn503,end_cn504,end_cn505,end_cn506,end_cn507,end_cn508,end_cn509,end_cn510,end_cn511,end_cn512,end_cn513,end_cn514,end_cn515,end_cn516,end_cn517,end_cn518,end_cn519,end_cn520,end_cn521,end_cn522,end_cn523,end_cn524,end_cn525,end_cn526,end_cn527,end_cn528,end_cn529,end_cn530,end_cn531,end_cn532,end_cn533,end_cn534,end_cn535,end_cn536,end_cn537,end_cn538,end_cn539,end_cn540,end_cn541,end_cn542,end_cn543,end_cn544,end_cn545,end_cn546,end_cn547,end_cn548,end_cn549,end_cn550,end_cn551,end_cn552,end_cn553,end_cn554,end_cn555,end_cn556,end_cn557,end_cn558,end_cn559,end_cn560,end_cn561,end_cn562,end_cn563,end_cn564,end_cn565,end_cn566,end_cn567,end_cn568,end_cn569,end_cn570,end_cn571,end_cn572,end_cn573,end_cn574,end_cn575,end_cn576,end_cn577,end_cn578,end_cn579,end_cn580,end_cn581,end_cn582,end_cn583,end_cn584,end_cn585,end_cn586,end_cn587,end_cn588,end_cn589,end_cn590,end_cn591,end_cn592,end_cn593,end_cn594,end_cn595,end_cn596,end_cn597,end_cn598,end_cn599,end_cn600,end_cn601,end_cn602,end_cn603,end_cn604,end_cn605,end_cn606,end_cn607,end_cn608,end_cn609,end_cn610,end_cn611,end_cn612,end_cn613,end_cn614,end_cn615,end_cn616,end_cn617,end_cn618,end_cn619,end_cn620,end_cn621,end_cn622,end_cn623,end_cn624,end_cn625,end_cn626,end_cn627,end_cn628,end_cn629,end_cn630,end_cn631,end_cn632,end_cn633,end_cn634,end_cn635,end_cn636,end_cn637,end_cn638,end_cn639,end_cn640,end_cn641,end_cn642,end_cn643,end_cn644,end_cn645,end_cn646,end_cn647,end_cn648,end_cn649,end_cn650,end_cn651,end_cn652,end_cn653,end_cn654,end_cn655,end_cn656,end_cn657,end_cn658,end_cn659,end_cn660,end_cn661,end_cn662,end_cn663,end_cn664,end_cn665,end_cn666,end_cn667,end_cn668,end_cn669,end_cn670,end_cn671,end_cn672,end_cn673,end_cn674,end_cn675,end_cn676,end_cn677,end_cn678,end_cn679,end_cn680,end_cn681,end_cn682,end_cn683,end_cn684,end_cn685,end_cn686,end_cn687,end_cn688,end_cn689,end_cn690,end_cn691,end_cn692,end_cn693,end_cn694,end_cn695,end_cn696,end_cn697,end_cn698,end_cn699,end_cn700,end_cn701,end_cn702,end_cn703,end_cn704,end_cn705,end_cn706,end_cn707,end_cn708,end_cn709,end_cn710,end_cn711,end_cn712,end_cn713,end_cn714,end_cn715,end_cn716,end_cn717,end_cn718,end_cn719,end_cn720,end_cn721,end_cn722,end_cn723,end_cn724,end_cn725,end_cn726,end_cn727,end_cn728,end_cn729,end_cn730,end_cn731,end_cn732,end_cn733,end_cn734,end_cn735,end_cn736,end_cn737,end_cn738,end_cn739,end_cn740,end_cn741,end_cn742,end_cn743,end_cn744,end_cn745,end_cn746,end_cn747,end_cn748,end_cn749,end_cn750,end_cn751,end_cn752,end_cn753,end_cn754,end_cn755,end_cn756,end_cn757,end_cn758,end_cn759,end_cn760,end_cn761,end_cn762,end_cn763,end_cn764,end_cn765,end_cn766,end_cn767,end_cn768,end_cn769,end_cn770,end_cn771,end_cn772,end_cn773,end_cn774,end_cn775,end_cn776,end_cn777,end_cn778,end_cn779,end_cn780,end_cn781,end_cn782,end_cn783,end_cn784,end_cn785,end_cn786,end_cn787,end_cn788,end_cn789,end_cn790,end_cn791,end_cn792,end_cn793,end_cn794,end_cn795,end_cn796,end_cn797,end_cn798,end_cn799,end_cn800,end_cn801,end_cn802,end_cn803,end_cn804,end_cn805,end_cn806,end_cn807,end_cn808,end_cn809,end_cn810,end_cn811,end_cn812,end_cn813,end_cn814,end_cn815,end_cn816,end_cn817,end_cn818,end_cn819,end_cn820,end_cn821,end_cn822,end_cn823,end_cn824,end_cn825,end_cn826,end_cn827,end_cn828,end_cn829,end_cn830,end_cn831,end_cn832,end_cn833,end_cn834,end_cn835,end_cn836,end_cn837,end_cn838,end_cn839,end_cn840,end_cn841,end_cn842,end_cn843,end_cn844,end_cn845,end_cn846,end_cn847,end_cn848,end_cn849,end_cn850,end_cn851,end_cn852,end_cn853,end_cn854,end_cn855,end_cn856,end_cn857,end_cn858,end_cn859,end_cn860,end_cn861,end_cn862,end_cn863,end_cn864,end_cn865,end_cn866,end_cn867,end_cn868,end_cn869,end_cn870,end_cn871,end_cn872,end_cn873,end_cn874,end_cn875,end_cn876,end_cn877,end_cn878,end_cn879,end_cn880,end_cn881,end_cn882,end_cn883,end_cn884,end_cn885,end_cn886,end_cn887,end_cn888,end_cn889,end_cn890,end_cn891,end_cn892,end_cn893,end_cn894,end_cn895,end_cn896,end_cn897,end_cn898,end_cn899,end_cn900,end_cn901,end_cn902,end_cn903,end_cn904,end_cn905,end_cn906,end_cn907,end_cn908,end_cn909,end_cn910,end_cn911,end_cn912,end_cn913,end_cn914,end_cn915,end_cn916,end_cn917,end_cn918,end_cn919,end_cn920,end_cn921,end_cn922,end_cn923,end_cn924,end_cn925,end_cn926,end_cn927,end_cn928,end_cn929,end_cn930,end_cn931,end_cn932,end_cn933,end_cn934,end_cn935,end_cn936,end_cn937,end_cn938,end_cn939,end_cn940,end_cn941,end_cn942,end_cn943,end_cn944,end_cn945,end_cn946,end_cn947,end_cn948,end_cn949,end_cn950,end_cn951,end_cn952,end_cn953,end_cn954,end_cn955,end_cn956,end_cn957,end_cn958,end_cn959,end_cn960,end_cn961,end_cn962,end_cn963,end_cn964,end_cn965,end_cn966,end_cn967,end_cn968,end_cn969,end_cn970,end_cn971,end_cn972,end_cn973,end_cn974,end_cn975,end_cn976,end_cn977,end_cn978,end_cn979,end_cn980,end_cn981,end_cn982,end_cn983,end_cn984,end_cn985,end_cn986,end_cn987,end_cn988,end_cn989,end_cn990,end_cn991,end_cn992,end_cn993,end_cn994,end_cn995,end_cn996,end_cn997,end_cn998,end_cn999,end_cn1000,end_cn1001,end_cn1002,end_cn1003,end_cn1004,end_cn1005,end_cn1006,end_cn1007,end_cn1008,end_cn1009,end_cn1010,end_cn1011,end_cn1012,end_cn1013,end_cn1014,end_cn1015,end_cn1016,end_cn1017,end_cn1018,end_cn1019,end_cn1020,end_cn1021,end_cn1022,end_cn1023,end_cn1024,end_cn1025,end_cn1026,end_cn1027,end_cn1028,end_cn1029,end_cn1030,end_cn1031,end_cn1032,end_cn1033,end_cn1034,end_cn1035,end_cn1036,end_cn1037,end_cn1038,end_cn1039,end_cn1040,end_cn1041,end_cn1042,end_cn1043,end_cn1044,end_cn1045,end_cn1046,end_cn1047,end_cn1048,end_cn1049,end_cn1050,end_cn1051,end_cn1052,end_cn1053,end_cn1054,end_cn1055,end_cn1056,end_cn1057,end_cn1058,end_cn1059,end_cn1060,end_cn1061,end_cn1062,end_cn1063,end_cn1064,end_cn1065,end_cn1066,end_cn1067,end_cn1068,end_cn1069,end_cn1070,end_cn1071,end_cn1072,end_cn1073,end_cn1074,end_cn1075,end_cn1076,end_cn1077,end_cn1078,end_cn1079,end_cn1080,end_cn1081,end_cn1082,end_cn1083,end_cn1084,end_cn1085,end_cn1086,end_cn1087,end_cn1088,end_cn1089,end_cn1090,end_cn1091,end_cn1092,end_cn1093,end_cn1094,end_cn1095,end_cn1096,end_cn1097,end_cn1098,end_cn1099,end_cn1100,end_cn1101,end_cn1102,end_cn1103,end_cn1104,end_cn1105,end_cn1106,end_cn1107,end_cn1108,end_cn1109,end_cn1110,end_cn1111,end_cn1112,end_cn1113,end_cn1114,end_cn1115,end_cn1116,end_cn1117,end_cn1118,end_cn1119,end_cn1120,end_cn1121,end_cn1122,end_cn1123,end_cn1124,end_cn1125,end_cn1126,end_cn1127,end_cn1128,end_cn1129,end_cn1130,end_cn1131,end_cn1132,end_cn1133,end_cn1134,end_cn1135,end_cn1136,end_cn1137,end_cn1138,end_cn1139,end_cn1140,end_cn1141,end_cn1142,end_cn1143,end_cn1144,end_cn1145,end_cn1146,end_cn1147,end_cn1148,end_cn1149,end_cn1150,end_cn1151,end_cn1152:std_logic;
begin
C1:CNPU6_6 port map (start_cn,clk,rst,V191C1,V266C1,V824C1,V948C1,V1160C1,V1249C1,C1V191,C1V266,C1V824,C1V948,C1V1160,C1V1249,end_cn1);
C2:CNPU6_6 port map (start_cn,clk,rst,V192C2,V267C2,V825C2,V949C2,V1161C2,V1250C2,C2V192,C2V267,C2V825,C2V949,C2V1161,C2V1250,end_cn2);
C3:CNPU6_6 port map (start_cn,clk,rst,V97C3,V268C3,V826C3,V950C3,V1162C3,V1251C3,C3V97,C3V268,C3V826,C3V950,C3V1162,C3V1251,end_cn3);
C4:CNPU6_6 port map (start_cn,clk,rst,V98C4,V269C4,V827C4,V951C4,V1163C4,V1252C4,C4V98,C4V269,C4V827,C4V951,C4V1163,C4V1252,end_cn4);
C5:CNPU6_6 port map (start_cn,clk,rst,V99C5,V270C5,V828C5,V952C5,V1164C5,V1253C5,C5V99,C5V270,C5V828,C5V952,C5V1164,C5V1253,end_cn5);
C6:CNPU6_6 port map (start_cn,clk,rst,V100C6,V271C6,V829C6,V953C6,V1165C6,V1254C6,C6V100,C6V271,C6V829,C6V953,C6V1165,C6V1254,end_cn6);
C7:CNPU6_6 port map (start_cn,clk,rst,V101C7,V272C7,V830C7,V954C7,V1166C7,V1255C7,C7V101,C7V272,C7V830,C7V954,C7V1166,C7V1255,end_cn7);
C8:CNPU6_6 port map (start_cn,clk,rst,V102C8,V273C8,V831C8,V955C8,V1167C8,V1256C8,C8V102,C8V273,C8V831,C8V955,C8V1167,C8V1256,end_cn8);
C9:CNPU6_6 port map (start_cn,clk,rst,V103C9,V274C9,V832C9,V956C9,V1168C9,V1257C9,C9V103,C9V274,C9V832,C9V956,C9V1168,C9V1257,end_cn9);
C10:CNPU6_6 port map (start_cn,clk,rst,V104C10,V275C10,V833C10,V957C10,V1169C10,V1258C10,C10V104,C10V275,C10V833,C10V957,C10V1169,C10V1258,end_cn10);
C11:CNPU6_6 port map (start_cn,clk,rst,V105C11,V276C11,V834C11,V958C11,V1170C11,V1259C11,C11V105,C11V276,C11V834,C11V958,C11V1170,C11V1259,end_cn11);
C12:CNPU6_6 port map (start_cn,clk,rst,V106C12,V277C12,V835C12,V959C12,V1171C12,V1260C12,C12V106,C12V277,C12V835,C12V959,C12V1171,C12V1260,end_cn12);
C13:CNPU6_6 port map (start_cn,clk,rst,V107C13,V278C13,V836C13,V960C13,V1172C13,V1261C13,C13V107,C13V278,C13V836,C13V960,C13V1172,C13V1261,end_cn13);
C14:CNPU6_6 port map (start_cn,clk,rst,V108C14,V279C14,V837C14,V865C14,V1173C14,V1262C14,C14V108,C14V279,C14V837,C14V865,C14V1173,C14V1262,end_cn14);
C15:CNPU6_6 port map (start_cn,clk,rst,V109C15,V280C15,V838C15,V866C15,V1174C15,V1263C15,C15V109,C15V280,C15V838,C15V866,C15V1174,C15V1263,end_cn15);
C16:CNPU6_6 port map (start_cn,clk,rst,V110C16,V281C16,V839C16,V867C16,V1175C16,V1264C16,C16V110,C16V281,C16V839,C16V867,C16V1175,C16V1264,end_cn16);
C17:CNPU6_6 port map (start_cn,clk,rst,V111C17,V282C17,V840C17,V868C17,V1176C17,V1265C17,C17V111,C17V282,C17V840,C17V868,C17V1176,C17V1265,end_cn17);
C18:CNPU6_6 port map (start_cn,clk,rst,V112C18,V283C18,V841C18,V869C18,V1177C18,V1266C18,C18V112,C18V283,C18V841,C18V869,C18V1177,C18V1266,end_cn18);
C19:CNPU6_6 port map (start_cn,clk,rst,V113C19,V284C19,V842C19,V870C19,V1178C19,V1267C19,C19V113,C19V284,C19V842,C19V870,C19V1178,C19V1267,end_cn19);
C20:CNPU6_6 port map (start_cn,clk,rst,V114C20,V285C20,V843C20,V871C20,V1179C20,V1268C20,C20V114,C20V285,C20V843,C20V871,C20V1179,C20V1268,end_cn20);
C21:CNPU6_6 port map (start_cn,clk,rst,V115C21,V286C21,V844C21,V872C21,V1180C21,V1269C21,C21V115,C21V286,C21V844,C21V872,C21V1180,C21V1269,end_cn21);
C22:CNPU6_6 port map (start_cn,clk,rst,V116C22,V287C22,V845C22,V873C22,V1181C22,V1270C22,C22V116,C22V287,C22V845,C22V873,C22V1181,C22V1270,end_cn22);
C23:CNPU6_6 port map (start_cn,clk,rst,V117C23,V288C23,V846C23,V874C23,V1182C23,V1271C23,C23V117,C23V288,C23V846,C23V874,C23V1182,C23V1271,end_cn23);
C24:CNPU6_6 port map (start_cn,clk,rst,V118C24,V193C24,V847C24,V875C24,V1183C24,V1272C24,C24V118,C24V193,C24V847,C24V875,C24V1183,C24V1272,end_cn24);
C25:CNPU6_6 port map (start_cn,clk,rst,V119C25,V194C25,V848C25,V876C25,V1184C25,V1273C25,C25V119,C25V194,C25V848,C25V876,C25V1184,C25V1273,end_cn25);
C26:CNPU6_6 port map (start_cn,clk,rst,V120C26,V195C26,V849C26,V877C26,V1185C26,V1274C26,C26V120,C26V195,C26V849,C26V877,C26V1185,C26V1274,end_cn26);
C27:CNPU6_6 port map (start_cn,clk,rst,V121C27,V196C27,V850C27,V878C27,V1186C27,V1275C27,C27V121,C27V196,C27V850,C27V878,C27V1186,C27V1275,end_cn27);
C28:CNPU6_6 port map (start_cn,clk,rst,V122C28,V197C28,V851C28,V879C28,V1187C28,V1276C28,C28V122,C28V197,C28V851,C28V879,C28V1187,C28V1276,end_cn28);
C29:CNPU6_6 port map (start_cn,clk,rst,V123C29,V198C29,V852C29,V880C29,V1188C29,V1277C29,C29V123,C29V198,C29V852,C29V880,C29V1188,C29V1277,end_cn29);
C30:CNPU6_6 port map (start_cn,clk,rst,V124C30,V199C30,V853C30,V881C30,V1189C30,V1278C30,C30V124,C30V199,C30V853,C30V881,C30V1189,C30V1278,end_cn30);
C31:CNPU6_6 port map (start_cn,clk,rst,V125C31,V200C31,V854C31,V882C31,V1190C31,V1279C31,C31V125,C31V200,C31V854,C31V882,C31V1190,C31V1279,end_cn31);
C32:CNPU6_6 port map (start_cn,clk,rst,V126C32,V201C32,V855C32,V883C32,V1191C32,V1280C32,C32V126,C32V201,C32V855,C32V883,C32V1191,C32V1280,end_cn32);
C33:CNPU6_6 port map (start_cn,clk,rst,V127C33,V202C33,V856C33,V884C33,V1192C33,V1281C33,C33V127,C33V202,C33V856,C33V884,C33V1192,C33V1281,end_cn33);
C34:CNPU6_6 port map (start_cn,clk,rst,V128C34,V203C34,V857C34,V885C34,V1193C34,V1282C34,C34V128,C34V203,C34V857,C34V885,C34V1193,C34V1282,end_cn34);
C35:CNPU6_6 port map (start_cn,clk,rst,V129C35,V204C35,V858C35,V886C35,V1194C35,V1283C35,C35V129,C35V204,C35V858,C35V886,C35V1194,C35V1283,end_cn35);
C36:CNPU6_6 port map (start_cn,clk,rst,V130C36,V205C36,V859C36,V887C36,V1195C36,V1284C36,C36V130,C36V205,C36V859,C36V887,C36V1195,C36V1284,end_cn36);
C37:CNPU6_6 port map (start_cn,clk,rst,V131C37,V206C37,V860C37,V888C37,V1196C37,V1285C37,C37V131,C37V206,C37V860,C37V888,C37V1196,C37V1285,end_cn37);
C38:CNPU6_6 port map (start_cn,clk,rst,V132C38,V207C38,V861C38,V889C38,V1197C38,V1286C38,C38V132,C38V207,C38V861,C38V889,C38V1197,C38V1286,end_cn38);
C39:CNPU6_6 port map (start_cn,clk,rst,V133C39,V208C39,V862C39,V890C39,V1198C39,V1287C39,C39V133,C39V208,C39V862,C39V890,C39V1198,C39V1287,end_cn39);
C40:CNPU6_6 port map (start_cn,clk,rst,V134C40,V209C40,V863C40,V891C40,V1199C40,V1288C40,C40V134,C40V209,C40V863,C40V891,C40V1199,C40V1288,end_cn40);
C41:CNPU6_6 port map (start_cn,clk,rst,V135C41,V210C41,V864C41,V892C41,V1200C41,V1289C41,C41V135,C41V210,C41V864,C41V892,C41V1200,C41V1289,end_cn41);
C42:CNPU6_6 port map (start_cn,clk,rst,V136C42,V211C42,V769C42,V893C42,V1201C42,V1290C42,C42V136,C42V211,C42V769,C42V893,C42V1201,C42V1290,end_cn42);
C43:CNPU6_6 port map (start_cn,clk,rst,V137C43,V212C43,V770C43,V894C43,V1202C43,V1291C43,C43V137,C43V212,C43V770,C43V894,C43V1202,C43V1291,end_cn43);
C44:CNPU6_6 port map (start_cn,clk,rst,V138C44,V213C44,V771C44,V895C44,V1203C44,V1292C44,C44V138,C44V213,C44V771,C44V895,C44V1203,C44V1292,end_cn44);
C45:CNPU6_6 port map (start_cn,clk,rst,V139C45,V214C45,V772C45,V896C45,V1204C45,V1293C45,C45V139,C45V214,C45V772,C45V896,C45V1204,C45V1293,end_cn45);
C46:CNPU6_6 port map (start_cn,clk,rst,V140C46,V215C46,V773C46,V897C46,V1205C46,V1294C46,C46V140,C46V215,C46V773,C46V897,C46V1205,C46V1294,end_cn46);
C47:CNPU6_6 port map (start_cn,clk,rst,V141C47,V216C47,V774C47,V898C47,V1206C47,V1295C47,C47V141,C47V216,C47V774,C47V898,C47V1206,C47V1295,end_cn47);
C48:CNPU6_6 port map (start_cn,clk,rst,V142C48,V217C48,V775C48,V899C48,V1207C48,V1296C48,C48V142,C48V217,C48V775,C48V899,C48V1207,C48V1296,end_cn48);
C49:CNPU6_6 port map (start_cn,clk,rst,V143C49,V218C49,V776C49,V900C49,V1208C49,V1297C49,C49V143,C49V218,C49V776,C49V900,C49V1208,C49V1297,end_cn49);
C50:CNPU6_6 port map (start_cn,clk,rst,V144C50,V219C50,V777C50,V901C50,V1209C50,V1298C50,C50V144,C50V219,C50V777,C50V901,C50V1209,C50V1298,end_cn50);
C51:CNPU6_6 port map (start_cn,clk,rst,V145C51,V220C51,V778C51,V902C51,V1210C51,V1299C51,C51V145,C51V220,C51V778,C51V902,C51V1210,C51V1299,end_cn51);
C52:CNPU6_6 port map (start_cn,clk,rst,V146C52,V221C52,V779C52,V903C52,V1211C52,V1300C52,C52V146,C52V221,C52V779,C52V903,C52V1211,C52V1300,end_cn52);
C53:CNPU6_6 port map (start_cn,clk,rst,V147C53,V222C53,V780C53,V904C53,V1212C53,V1301C53,C53V147,C53V222,C53V780,C53V904,C53V1212,C53V1301,end_cn53);
C54:CNPU6_6 port map (start_cn,clk,rst,V148C54,V223C54,V781C54,V905C54,V1213C54,V1302C54,C54V148,C54V223,C54V781,C54V905,C54V1213,C54V1302,end_cn54);
C55:CNPU6_6 port map (start_cn,clk,rst,V149C55,V224C55,V782C55,V906C55,V1214C55,V1303C55,C55V149,C55V224,C55V782,C55V906,C55V1214,C55V1303,end_cn55);
C56:CNPU6_6 port map (start_cn,clk,rst,V150C56,V225C56,V783C56,V907C56,V1215C56,V1304C56,C56V150,C56V225,C56V783,C56V907,C56V1215,C56V1304,end_cn56);
C57:CNPU6_6 port map (start_cn,clk,rst,V151C57,V226C57,V784C57,V908C57,V1216C57,V1305C57,C57V151,C57V226,C57V784,C57V908,C57V1216,C57V1305,end_cn57);
C58:CNPU6_6 port map (start_cn,clk,rst,V152C58,V227C58,V785C58,V909C58,V1217C58,V1306C58,C58V152,C58V227,C58V785,C58V909,C58V1217,C58V1306,end_cn58);
C59:CNPU6_6 port map (start_cn,clk,rst,V153C59,V228C59,V786C59,V910C59,V1218C59,V1307C59,C59V153,C59V228,C59V786,C59V910,C59V1218,C59V1307,end_cn59);
C60:CNPU6_6 port map (start_cn,clk,rst,V154C60,V229C60,V787C60,V911C60,V1219C60,V1308C60,C60V154,C60V229,C60V787,C60V911,C60V1219,C60V1308,end_cn60);
C61:CNPU6_6 port map (start_cn,clk,rst,V155C61,V230C61,V788C61,V912C61,V1220C61,V1309C61,C61V155,C61V230,C61V788,C61V912,C61V1220,C61V1309,end_cn61);
C62:CNPU6_6 port map (start_cn,clk,rst,V156C62,V231C62,V789C62,V913C62,V1221C62,V1310C62,C62V156,C62V231,C62V789,C62V913,C62V1221,C62V1310,end_cn62);
C63:CNPU6_6 port map (start_cn,clk,rst,V157C63,V232C63,V790C63,V914C63,V1222C63,V1311C63,C63V157,C63V232,C63V790,C63V914,C63V1222,C63V1311,end_cn63);
C64:CNPU6_6 port map (start_cn,clk,rst,V158C64,V233C64,V791C64,V915C64,V1223C64,V1312C64,C64V158,C64V233,C64V791,C64V915,C64V1223,C64V1312,end_cn64);
C65:CNPU6_6 port map (start_cn,clk,rst,V159C65,V234C65,V792C65,V916C65,V1224C65,V1313C65,C65V159,C65V234,C65V792,C65V916,C65V1224,C65V1313,end_cn65);
C66:CNPU6_6 port map (start_cn,clk,rst,V160C66,V235C66,V793C66,V917C66,V1225C66,V1314C66,C66V160,C66V235,C66V793,C66V917,C66V1225,C66V1314,end_cn66);
C67:CNPU6_6 port map (start_cn,clk,rst,V161C67,V236C67,V794C67,V918C67,V1226C67,V1315C67,C67V161,C67V236,C67V794,C67V918,C67V1226,C67V1315,end_cn67);
C68:CNPU6_6 port map (start_cn,clk,rst,V162C68,V237C68,V795C68,V919C68,V1227C68,V1316C68,C68V162,C68V237,C68V795,C68V919,C68V1227,C68V1316,end_cn68);
C69:CNPU6_6 port map (start_cn,clk,rst,V163C69,V238C69,V796C69,V920C69,V1228C69,V1317C69,C69V163,C69V238,C69V796,C69V920,C69V1228,C69V1317,end_cn69);
C70:CNPU6_6 port map (start_cn,clk,rst,V164C70,V239C70,V797C70,V921C70,V1229C70,V1318C70,C70V164,C70V239,C70V797,C70V921,C70V1229,C70V1318,end_cn70);
C71:CNPU6_6 port map (start_cn,clk,rst,V165C71,V240C71,V798C71,V922C71,V1230C71,V1319C71,C71V165,C71V240,C71V798,C71V922,C71V1230,C71V1319,end_cn71);
C72:CNPU6_6 port map (start_cn,clk,rst,V166C72,V241C72,V799C72,V923C72,V1231C72,V1320C72,C72V166,C72V241,C72V799,C72V923,C72V1231,C72V1320,end_cn72);
C73:CNPU6_6 port map (start_cn,clk,rst,V167C73,V242C73,V800C73,V924C73,V1232C73,V1321C73,C73V167,C73V242,C73V800,C73V924,C73V1232,C73V1321,end_cn73);
C74:CNPU6_6 port map (start_cn,clk,rst,V168C74,V243C74,V801C74,V925C74,V1233C74,V1322C74,C74V168,C74V243,C74V801,C74V925,C74V1233,C74V1322,end_cn74);
C75:CNPU6_6 port map (start_cn,clk,rst,V169C75,V244C75,V802C75,V926C75,V1234C75,V1323C75,C75V169,C75V244,C75V802,C75V926,C75V1234,C75V1323,end_cn75);
C76:CNPU6_6 port map (start_cn,clk,rst,V170C76,V245C76,V803C76,V927C76,V1235C76,V1324C76,C76V170,C76V245,C76V803,C76V927,C76V1235,C76V1324,end_cn76);
C77:CNPU6_6 port map (start_cn,clk,rst,V171C77,V246C77,V804C77,V928C77,V1236C77,V1325C77,C77V171,C77V246,C77V804,C77V928,C77V1236,C77V1325,end_cn77);
C78:CNPU6_6 port map (start_cn,clk,rst,V172C78,V247C78,V805C78,V929C78,V1237C78,V1326C78,C78V172,C78V247,C78V805,C78V929,C78V1237,C78V1326,end_cn78);
C79:CNPU6_6 port map (start_cn,clk,rst,V173C79,V248C79,V806C79,V930C79,V1238C79,V1327C79,C79V173,C79V248,C79V806,C79V930,C79V1238,C79V1327,end_cn79);
C80:CNPU6_6 port map (start_cn,clk,rst,V174C80,V249C80,V807C80,V931C80,V1239C80,V1328C80,C80V174,C80V249,C80V807,C80V931,C80V1239,C80V1328,end_cn80);
C81:CNPU6_6 port map (start_cn,clk,rst,V175C81,V250C81,V808C81,V932C81,V1240C81,V1329C81,C81V175,C81V250,C81V808,C81V932,C81V1240,C81V1329,end_cn81);
C82:CNPU6_6 port map (start_cn,clk,rst,V176C82,V251C82,V809C82,V933C82,V1241C82,V1330C82,C82V176,C82V251,C82V809,C82V933,C82V1241,C82V1330,end_cn82);
C83:CNPU6_6 port map (start_cn,clk,rst,V177C83,V252C83,V810C83,V934C83,V1242C83,V1331C83,C83V177,C83V252,C83V810,C83V934,C83V1242,C83V1331,end_cn83);
C84:CNPU6_6 port map (start_cn,clk,rst,V178C84,V253C84,V811C84,V935C84,V1243C84,V1332C84,C84V178,C84V253,C84V811,C84V935,C84V1243,C84V1332,end_cn84);
C85:CNPU6_6 port map (start_cn,clk,rst,V179C85,V254C85,V812C85,V936C85,V1244C85,V1333C85,C85V179,C85V254,C85V812,C85V936,C85V1244,C85V1333,end_cn85);
C86:CNPU6_6 port map (start_cn,clk,rst,V180C86,V255C86,V813C86,V937C86,V1245C86,V1334C86,C86V180,C86V255,C86V813,C86V937,C86V1245,C86V1334,end_cn86);
C87:CNPU6_6 port map (start_cn,clk,rst,V181C87,V256C87,V814C87,V938C87,V1246C87,V1335C87,C87V181,C87V256,C87V814,C87V938,C87V1246,C87V1335,end_cn87);
C88:CNPU6_6 port map (start_cn,clk,rst,V182C88,V257C88,V815C88,V939C88,V1247C88,V1336C88,C88V182,C88V257,C88V815,C88V939,C88V1247,C88V1336,end_cn88);
C89:CNPU6_6 port map (start_cn,clk,rst,V183C89,V258C89,V816C89,V940C89,V1248C89,V1337C89,C89V183,C89V258,C89V816,C89V940,C89V1248,C89V1337,end_cn89);
C90:CNPU6_6 port map (start_cn,clk,rst,V184C90,V259C90,V817C90,V941C90,V1153C90,V1338C90,C90V184,C90V259,C90V817,C90V941,C90V1153,C90V1338,end_cn90);
C91:CNPU6_6 port map (start_cn,clk,rst,V185C91,V260C91,V818C91,V942C91,V1154C91,V1339C91,C91V185,C91V260,C91V818,C91V942,C91V1154,C91V1339,end_cn91);
C92:CNPU6_6 port map (start_cn,clk,rst,V186C92,V261C92,V819C92,V943C92,V1155C92,V1340C92,C92V186,C92V261,C92V819,C92V943,C92V1155,C92V1340,end_cn92);
C93:CNPU6_6 port map (start_cn,clk,rst,V187C93,V262C93,V820C93,V944C93,V1156C93,V1341C93,C93V187,C93V262,C93V820,C93V944,C93V1156,C93V1341,end_cn93);
C94:CNPU6_6 port map (start_cn,clk,rst,V188C94,V263C94,V821C94,V945C94,V1157C94,V1342C94,C94V188,C94V263,C94V821,C94V945,C94V1157,C94V1342,end_cn94);
C95:CNPU6_6 port map (start_cn,clk,rst,V189C95,V264C95,V822C95,V946C95,V1158C95,V1343C95,C95V189,C95V264,C95V822,C95V946,C95V1158,C95V1343,end_cn95);
C96:CNPU6_6 port map (start_cn,clk,rst,V190C96,V265C96,V823C96,V947C96,V1159C96,V1344C96,C96V190,C96V265,C96V823,C96V947,C96V1159,C96V1344,end_cn96);
C97:CNPU7_7 port map (start_cn,clk,rst,V124C97,V503C97,V656C97,V682C97,V1069C97,V1249C97,V1345C97,C97V124,C97V503,C97V656,C97V682,C97V1069,C97V1249,C97V1345,end_cn97);
C98:CNPU7_7 port map (start_cn,clk,rst,V125C98,V504C98,V657C98,V683C98,V1070C98,V1250C98,V1346C98,C98V125,C98V504,C98V657,C98V683,C98V1070,C98V1250,C98V1346,end_cn98);
C99:CNPU7_7 port map (start_cn,clk,rst,V126C99,V505C99,V658C99,V684C99,V1071C99,V1251C99,V1347C99,C99V126,C99V505,C99V658,C99V684,C99V1071,C99V1251,C99V1347,end_cn99);
C100:CNPU7_7 port map (start_cn,clk,rst,V127C100,V506C100,V659C100,V685C100,V1072C100,V1252C100,V1348C100,C100V127,C100V506,C100V659,C100V685,C100V1072,C100V1252,C100V1348,end_cn100);
C101:CNPU7_7 port map (start_cn,clk,rst,V128C101,V507C101,V660C101,V686C101,V1073C101,V1253C101,V1349C101,C101V128,C101V507,C101V660,C101V686,C101V1073,C101V1253,C101V1349,end_cn101);
C102:CNPU7_7 port map (start_cn,clk,rst,V129C102,V508C102,V661C102,V687C102,V1074C102,V1254C102,V1350C102,C102V129,C102V508,C102V661,C102V687,C102V1074,C102V1254,C102V1350,end_cn102);
C103:CNPU7_7 port map (start_cn,clk,rst,V130C103,V509C103,V662C103,V688C103,V1075C103,V1255C103,V1351C103,C103V130,C103V509,C103V662,C103V688,C103V1075,C103V1255,C103V1351,end_cn103);
C104:CNPU7_7 port map (start_cn,clk,rst,V131C104,V510C104,V663C104,V689C104,V1076C104,V1256C104,V1352C104,C104V131,C104V510,C104V663,C104V689,C104V1076,C104V1256,C104V1352,end_cn104);
C105:CNPU7_7 port map (start_cn,clk,rst,V132C105,V511C105,V664C105,V690C105,V1077C105,V1257C105,V1353C105,C105V132,C105V511,C105V664,C105V690,C105V1077,C105V1257,C105V1353,end_cn105);
C106:CNPU7_7 port map (start_cn,clk,rst,V133C106,V512C106,V665C106,V691C106,V1078C106,V1258C106,V1354C106,C106V133,C106V512,C106V665,C106V691,C106V1078,C106V1258,C106V1354,end_cn106);
C107:CNPU7_7 port map (start_cn,clk,rst,V134C107,V513C107,V666C107,V692C107,V1079C107,V1259C107,V1355C107,C107V134,C107V513,C107V666,C107V692,C107V1079,C107V1259,C107V1355,end_cn107);
C108:CNPU7_7 port map (start_cn,clk,rst,V135C108,V514C108,V667C108,V693C108,V1080C108,V1260C108,V1356C108,C108V135,C108V514,C108V667,C108V693,C108V1080,C108V1260,C108V1356,end_cn108);
C109:CNPU7_7 port map (start_cn,clk,rst,V136C109,V515C109,V668C109,V694C109,V1081C109,V1261C109,V1357C109,C109V136,C109V515,C109V668,C109V694,C109V1081,C109V1261,C109V1357,end_cn109);
C110:CNPU7_7 port map (start_cn,clk,rst,V137C110,V516C110,V669C110,V695C110,V1082C110,V1262C110,V1358C110,C110V137,C110V516,C110V669,C110V695,C110V1082,C110V1262,C110V1358,end_cn110);
C111:CNPU7_7 port map (start_cn,clk,rst,V138C111,V517C111,V670C111,V696C111,V1083C111,V1263C111,V1359C111,C111V138,C111V517,C111V670,C111V696,C111V1083,C111V1263,C111V1359,end_cn111);
C112:CNPU7_7 port map (start_cn,clk,rst,V139C112,V518C112,V671C112,V697C112,V1084C112,V1264C112,V1360C112,C112V139,C112V518,C112V671,C112V697,C112V1084,C112V1264,C112V1360,end_cn112);
C113:CNPU7_7 port map (start_cn,clk,rst,V140C113,V519C113,V672C113,V698C113,V1085C113,V1265C113,V1361C113,C113V140,C113V519,C113V672,C113V698,C113V1085,C113V1265,C113V1361,end_cn113);
C114:CNPU7_7 port map (start_cn,clk,rst,V141C114,V520C114,V577C114,V699C114,V1086C114,V1266C114,V1362C114,C114V141,C114V520,C114V577,C114V699,C114V1086,C114V1266,C114V1362,end_cn114);
C115:CNPU7_7 port map (start_cn,clk,rst,V142C115,V521C115,V578C115,V700C115,V1087C115,V1267C115,V1363C115,C115V142,C115V521,C115V578,C115V700,C115V1087,C115V1267,C115V1363,end_cn115);
C116:CNPU7_7 port map (start_cn,clk,rst,V143C116,V522C116,V579C116,V701C116,V1088C116,V1268C116,V1364C116,C116V143,C116V522,C116V579,C116V701,C116V1088,C116V1268,C116V1364,end_cn116);
C117:CNPU7_7 port map (start_cn,clk,rst,V144C117,V523C117,V580C117,V702C117,V1089C117,V1269C117,V1365C117,C117V144,C117V523,C117V580,C117V702,C117V1089,C117V1269,C117V1365,end_cn117);
C118:CNPU7_7 port map (start_cn,clk,rst,V145C118,V524C118,V581C118,V703C118,V1090C118,V1270C118,V1366C118,C118V145,C118V524,C118V581,C118V703,C118V1090,C118V1270,C118V1366,end_cn118);
C119:CNPU7_7 port map (start_cn,clk,rst,V146C119,V525C119,V582C119,V704C119,V1091C119,V1271C119,V1367C119,C119V146,C119V525,C119V582,C119V704,C119V1091,C119V1271,C119V1367,end_cn119);
C120:CNPU7_7 port map (start_cn,clk,rst,V147C120,V526C120,V583C120,V705C120,V1092C120,V1272C120,V1368C120,C120V147,C120V526,C120V583,C120V705,C120V1092,C120V1272,C120V1368,end_cn120);
C121:CNPU7_7 port map (start_cn,clk,rst,V148C121,V527C121,V584C121,V706C121,V1093C121,V1273C121,V1369C121,C121V148,C121V527,C121V584,C121V706,C121V1093,C121V1273,C121V1369,end_cn121);
C122:CNPU7_7 port map (start_cn,clk,rst,V149C122,V528C122,V585C122,V707C122,V1094C122,V1274C122,V1370C122,C122V149,C122V528,C122V585,C122V707,C122V1094,C122V1274,C122V1370,end_cn122);
C123:CNPU7_7 port map (start_cn,clk,rst,V150C123,V529C123,V586C123,V708C123,V1095C123,V1275C123,V1371C123,C123V150,C123V529,C123V586,C123V708,C123V1095,C123V1275,C123V1371,end_cn123);
C124:CNPU7_7 port map (start_cn,clk,rst,V151C124,V530C124,V587C124,V709C124,V1096C124,V1276C124,V1372C124,C124V151,C124V530,C124V587,C124V709,C124V1096,C124V1276,C124V1372,end_cn124);
C125:CNPU7_7 port map (start_cn,clk,rst,V152C125,V531C125,V588C125,V710C125,V1097C125,V1277C125,V1373C125,C125V152,C125V531,C125V588,C125V710,C125V1097,C125V1277,C125V1373,end_cn125);
C126:CNPU7_7 port map (start_cn,clk,rst,V153C126,V532C126,V589C126,V711C126,V1098C126,V1278C126,V1374C126,C126V153,C126V532,C126V589,C126V711,C126V1098,C126V1278,C126V1374,end_cn126);
C127:CNPU7_7 port map (start_cn,clk,rst,V154C127,V533C127,V590C127,V712C127,V1099C127,V1279C127,V1375C127,C127V154,C127V533,C127V590,C127V712,C127V1099,C127V1279,C127V1375,end_cn127);
C128:CNPU7_7 port map (start_cn,clk,rst,V155C128,V534C128,V591C128,V713C128,V1100C128,V1280C128,V1376C128,C128V155,C128V534,C128V591,C128V713,C128V1100,C128V1280,C128V1376,end_cn128);
C129:CNPU7_7 port map (start_cn,clk,rst,V156C129,V535C129,V592C129,V714C129,V1101C129,V1281C129,V1377C129,C129V156,C129V535,C129V592,C129V714,C129V1101,C129V1281,C129V1377,end_cn129);
C130:CNPU7_7 port map (start_cn,clk,rst,V157C130,V536C130,V593C130,V715C130,V1102C130,V1282C130,V1378C130,C130V157,C130V536,C130V593,C130V715,C130V1102,C130V1282,C130V1378,end_cn130);
C131:CNPU7_7 port map (start_cn,clk,rst,V158C131,V537C131,V594C131,V716C131,V1103C131,V1283C131,V1379C131,C131V158,C131V537,C131V594,C131V716,C131V1103,C131V1283,C131V1379,end_cn131);
C132:CNPU7_7 port map (start_cn,clk,rst,V159C132,V538C132,V595C132,V717C132,V1104C132,V1284C132,V1380C132,C132V159,C132V538,C132V595,C132V717,C132V1104,C132V1284,C132V1380,end_cn132);
C133:CNPU7_7 port map (start_cn,clk,rst,V160C133,V539C133,V596C133,V718C133,V1105C133,V1285C133,V1381C133,C133V160,C133V539,C133V596,C133V718,C133V1105,C133V1285,C133V1381,end_cn133);
C134:CNPU7_7 port map (start_cn,clk,rst,V161C134,V540C134,V597C134,V719C134,V1106C134,V1286C134,V1382C134,C134V161,C134V540,C134V597,C134V719,C134V1106,C134V1286,C134V1382,end_cn134);
C135:CNPU7_7 port map (start_cn,clk,rst,V162C135,V541C135,V598C135,V720C135,V1107C135,V1287C135,V1383C135,C135V162,C135V541,C135V598,C135V720,C135V1107,C135V1287,C135V1383,end_cn135);
C136:CNPU7_7 port map (start_cn,clk,rst,V163C136,V542C136,V599C136,V721C136,V1108C136,V1288C136,V1384C136,C136V163,C136V542,C136V599,C136V721,C136V1108,C136V1288,C136V1384,end_cn136);
C137:CNPU7_7 port map (start_cn,clk,rst,V164C137,V543C137,V600C137,V722C137,V1109C137,V1289C137,V1385C137,C137V164,C137V543,C137V600,C137V722,C137V1109,C137V1289,C137V1385,end_cn137);
C138:CNPU7_7 port map (start_cn,clk,rst,V165C138,V544C138,V601C138,V723C138,V1110C138,V1290C138,V1386C138,C138V165,C138V544,C138V601,C138V723,C138V1110,C138V1290,C138V1386,end_cn138);
C139:CNPU7_7 port map (start_cn,clk,rst,V166C139,V545C139,V602C139,V724C139,V1111C139,V1291C139,V1387C139,C139V166,C139V545,C139V602,C139V724,C139V1111,C139V1291,C139V1387,end_cn139);
C140:CNPU7_7 port map (start_cn,clk,rst,V167C140,V546C140,V603C140,V725C140,V1112C140,V1292C140,V1388C140,C140V167,C140V546,C140V603,C140V725,C140V1112,C140V1292,C140V1388,end_cn140);
C141:CNPU7_7 port map (start_cn,clk,rst,V168C141,V547C141,V604C141,V726C141,V1113C141,V1293C141,V1389C141,C141V168,C141V547,C141V604,C141V726,C141V1113,C141V1293,C141V1389,end_cn141);
C142:CNPU7_7 port map (start_cn,clk,rst,V169C142,V548C142,V605C142,V727C142,V1114C142,V1294C142,V1390C142,C142V169,C142V548,C142V605,C142V727,C142V1114,C142V1294,C142V1390,end_cn142);
C143:CNPU7_7 port map (start_cn,clk,rst,V170C143,V549C143,V606C143,V728C143,V1115C143,V1295C143,V1391C143,C143V170,C143V549,C143V606,C143V728,C143V1115,C143V1295,C143V1391,end_cn143);
C144:CNPU7_7 port map (start_cn,clk,rst,V171C144,V550C144,V607C144,V729C144,V1116C144,V1296C144,V1392C144,C144V171,C144V550,C144V607,C144V729,C144V1116,C144V1296,C144V1392,end_cn144);
C145:CNPU7_7 port map (start_cn,clk,rst,V172C145,V551C145,V608C145,V730C145,V1117C145,V1297C145,V1393C145,C145V172,C145V551,C145V608,C145V730,C145V1117,C145V1297,C145V1393,end_cn145);
C146:CNPU7_7 port map (start_cn,clk,rst,V173C146,V552C146,V609C146,V731C146,V1118C146,V1298C146,V1394C146,C146V173,C146V552,C146V609,C146V731,C146V1118,C146V1298,C146V1394,end_cn146);
C147:CNPU7_7 port map (start_cn,clk,rst,V174C147,V553C147,V610C147,V732C147,V1119C147,V1299C147,V1395C147,C147V174,C147V553,C147V610,C147V732,C147V1119,C147V1299,C147V1395,end_cn147);
C148:CNPU7_7 port map (start_cn,clk,rst,V175C148,V554C148,V611C148,V733C148,V1120C148,V1300C148,V1396C148,C148V175,C148V554,C148V611,C148V733,C148V1120,C148V1300,C148V1396,end_cn148);
C149:CNPU7_7 port map (start_cn,clk,rst,V176C149,V555C149,V612C149,V734C149,V1121C149,V1301C149,V1397C149,C149V176,C149V555,C149V612,C149V734,C149V1121,C149V1301,C149V1397,end_cn149);
C150:CNPU7_7 port map (start_cn,clk,rst,V177C150,V556C150,V613C150,V735C150,V1122C150,V1302C150,V1398C150,C150V177,C150V556,C150V613,C150V735,C150V1122,C150V1302,C150V1398,end_cn150);
C151:CNPU7_7 port map (start_cn,clk,rst,V178C151,V557C151,V614C151,V736C151,V1123C151,V1303C151,V1399C151,C151V178,C151V557,C151V614,C151V736,C151V1123,C151V1303,C151V1399,end_cn151);
C152:CNPU7_7 port map (start_cn,clk,rst,V179C152,V558C152,V615C152,V737C152,V1124C152,V1304C152,V1400C152,C152V179,C152V558,C152V615,C152V737,C152V1124,C152V1304,C152V1400,end_cn152);
C153:CNPU7_7 port map (start_cn,clk,rst,V180C153,V559C153,V616C153,V738C153,V1125C153,V1305C153,V1401C153,C153V180,C153V559,C153V616,C153V738,C153V1125,C153V1305,C153V1401,end_cn153);
C154:CNPU7_7 port map (start_cn,clk,rst,V181C154,V560C154,V617C154,V739C154,V1126C154,V1306C154,V1402C154,C154V181,C154V560,C154V617,C154V739,C154V1126,C154V1306,C154V1402,end_cn154);
C155:CNPU7_7 port map (start_cn,clk,rst,V182C155,V561C155,V618C155,V740C155,V1127C155,V1307C155,V1403C155,C155V182,C155V561,C155V618,C155V740,C155V1127,C155V1307,C155V1403,end_cn155);
C156:CNPU7_7 port map (start_cn,clk,rst,V183C156,V562C156,V619C156,V741C156,V1128C156,V1308C156,V1404C156,C156V183,C156V562,C156V619,C156V741,C156V1128,C156V1308,C156V1404,end_cn156);
C157:CNPU7_7 port map (start_cn,clk,rst,V184C157,V563C157,V620C157,V742C157,V1129C157,V1309C157,V1405C157,C157V184,C157V563,C157V620,C157V742,C157V1129,C157V1309,C157V1405,end_cn157);
C158:CNPU7_7 port map (start_cn,clk,rst,V185C158,V564C158,V621C158,V743C158,V1130C158,V1310C158,V1406C158,C158V185,C158V564,C158V621,C158V743,C158V1130,C158V1310,C158V1406,end_cn158);
C159:CNPU7_7 port map (start_cn,clk,rst,V186C159,V565C159,V622C159,V744C159,V1131C159,V1311C159,V1407C159,C159V186,C159V565,C159V622,C159V744,C159V1131,C159V1311,C159V1407,end_cn159);
C160:CNPU7_7 port map (start_cn,clk,rst,V187C160,V566C160,V623C160,V745C160,V1132C160,V1312C160,V1408C160,C160V187,C160V566,C160V623,C160V745,C160V1132,C160V1312,C160V1408,end_cn160);
C161:CNPU7_7 port map (start_cn,clk,rst,V188C161,V567C161,V624C161,V746C161,V1133C161,V1313C161,V1409C161,C161V188,C161V567,C161V624,C161V746,C161V1133,C161V1313,C161V1409,end_cn161);
C162:CNPU7_7 port map (start_cn,clk,rst,V189C162,V568C162,V625C162,V747C162,V1134C162,V1314C162,V1410C162,C162V189,C162V568,C162V625,C162V747,C162V1134,C162V1314,C162V1410,end_cn162);
C163:CNPU7_7 port map (start_cn,clk,rst,V190C163,V569C163,V626C163,V748C163,V1135C163,V1315C163,V1411C163,C163V190,C163V569,C163V626,C163V748,C163V1135,C163V1315,C163V1411,end_cn163);
C164:CNPU7_7 port map (start_cn,clk,rst,V191C164,V570C164,V627C164,V749C164,V1136C164,V1316C164,V1412C164,C164V191,C164V570,C164V627,C164V749,C164V1136,C164V1316,C164V1412,end_cn164);
C165:CNPU7_7 port map (start_cn,clk,rst,V192C165,V571C165,V628C165,V750C165,V1137C165,V1317C165,V1413C165,C165V192,C165V571,C165V628,C165V750,C165V1137,C165V1317,C165V1413,end_cn165);
C166:CNPU7_7 port map (start_cn,clk,rst,V97C166,V572C166,V629C166,V751C166,V1138C166,V1318C166,V1414C166,C166V97,C166V572,C166V629,C166V751,C166V1138,C166V1318,C166V1414,end_cn166);
C167:CNPU7_7 port map (start_cn,clk,rst,V98C167,V573C167,V630C167,V752C167,V1139C167,V1319C167,V1415C167,C167V98,C167V573,C167V630,C167V752,C167V1139,C167V1319,C167V1415,end_cn167);
C168:CNPU7_7 port map (start_cn,clk,rst,V99C168,V574C168,V631C168,V753C168,V1140C168,V1320C168,V1416C168,C168V99,C168V574,C168V631,C168V753,C168V1140,C168V1320,C168V1416,end_cn168);
C169:CNPU7_7 port map (start_cn,clk,rst,V100C169,V575C169,V632C169,V754C169,V1141C169,V1321C169,V1417C169,C169V100,C169V575,C169V632,C169V754,C169V1141,C169V1321,C169V1417,end_cn169);
C170:CNPU7_7 port map (start_cn,clk,rst,V101C170,V576C170,V633C170,V755C170,V1142C170,V1322C170,V1418C170,C170V101,C170V576,C170V633,C170V755,C170V1142,C170V1322,C170V1418,end_cn170);
C171:CNPU7_7 port map (start_cn,clk,rst,V102C171,V481C171,V634C171,V756C171,V1143C171,V1323C171,V1419C171,C171V102,C171V481,C171V634,C171V756,C171V1143,C171V1323,C171V1419,end_cn171);
C172:CNPU7_7 port map (start_cn,clk,rst,V103C172,V482C172,V635C172,V757C172,V1144C172,V1324C172,V1420C172,C172V103,C172V482,C172V635,C172V757,C172V1144,C172V1324,C172V1420,end_cn172);
C173:CNPU7_7 port map (start_cn,clk,rst,V104C173,V483C173,V636C173,V758C173,V1145C173,V1325C173,V1421C173,C173V104,C173V483,C173V636,C173V758,C173V1145,C173V1325,C173V1421,end_cn173);
C174:CNPU7_7 port map (start_cn,clk,rst,V105C174,V484C174,V637C174,V759C174,V1146C174,V1326C174,V1422C174,C174V105,C174V484,C174V637,C174V759,C174V1146,C174V1326,C174V1422,end_cn174);
C175:CNPU7_7 port map (start_cn,clk,rst,V106C175,V485C175,V638C175,V760C175,V1147C175,V1327C175,V1423C175,C175V106,C175V485,C175V638,C175V760,C175V1147,C175V1327,C175V1423,end_cn175);
C176:CNPU7_7 port map (start_cn,clk,rst,V107C176,V486C176,V639C176,V761C176,V1148C176,V1328C176,V1424C176,C176V107,C176V486,C176V639,C176V761,C176V1148,C176V1328,C176V1424,end_cn176);
C177:CNPU7_7 port map (start_cn,clk,rst,V108C177,V487C177,V640C177,V762C177,V1149C177,V1329C177,V1425C177,C177V108,C177V487,C177V640,C177V762,C177V1149,C177V1329,C177V1425,end_cn177);
C178:CNPU7_7 port map (start_cn,clk,rst,V109C178,V488C178,V641C178,V763C178,V1150C178,V1330C178,V1426C178,C178V109,C178V488,C178V641,C178V763,C178V1150,C178V1330,C178V1426,end_cn178);
C179:CNPU7_7 port map (start_cn,clk,rst,V110C179,V489C179,V642C179,V764C179,V1151C179,V1331C179,V1427C179,C179V110,C179V489,C179V642,C179V764,C179V1151,C179V1331,C179V1427,end_cn179);
C180:CNPU7_7 port map (start_cn,clk,rst,V111C180,V490C180,V643C180,V765C180,V1152C180,V1332C180,V1428C180,C180V111,C180V490,C180V643,C180V765,C180V1152,C180V1332,C180V1428,end_cn180);
C181:CNPU7_7 port map (start_cn,clk,rst,V112C181,V491C181,V644C181,V766C181,V1057C181,V1333C181,V1429C181,C181V112,C181V491,C181V644,C181V766,C181V1057,C181V1333,C181V1429,end_cn181);
C182:CNPU7_7 port map (start_cn,clk,rst,V113C182,V492C182,V645C182,V767C182,V1058C182,V1334C182,V1430C182,C182V113,C182V492,C182V645,C182V767,C182V1058,C182V1334,C182V1430,end_cn182);
C183:CNPU7_7 port map (start_cn,clk,rst,V114C183,V493C183,V646C183,V768C183,V1059C183,V1335C183,V1431C183,C183V114,C183V493,C183V646,C183V768,C183V1059,C183V1335,C183V1431,end_cn183);
C184:CNPU7_7 port map (start_cn,clk,rst,V115C184,V494C184,V647C184,V673C184,V1060C184,V1336C184,V1432C184,C184V115,C184V494,C184V647,C184V673,C184V1060,C184V1336,C184V1432,end_cn184);
C185:CNPU7_7 port map (start_cn,clk,rst,V116C185,V495C185,V648C185,V674C185,V1061C185,V1337C185,V1433C185,C185V116,C185V495,C185V648,C185V674,C185V1061,C185V1337,C185V1433,end_cn185);
C186:CNPU7_7 port map (start_cn,clk,rst,V117C186,V496C186,V649C186,V675C186,V1062C186,V1338C186,V1434C186,C186V117,C186V496,C186V649,C186V675,C186V1062,C186V1338,C186V1434,end_cn186);
C187:CNPU7_7 port map (start_cn,clk,rst,V118C187,V497C187,V650C187,V676C187,V1063C187,V1339C187,V1435C187,C187V118,C187V497,C187V650,C187V676,C187V1063,C187V1339,C187V1435,end_cn187);
C188:CNPU7_7 port map (start_cn,clk,rst,V119C188,V498C188,V651C188,V677C188,V1064C188,V1340C188,V1436C188,C188V119,C188V498,C188V651,C188V677,C188V1064,C188V1340,C188V1436,end_cn188);
C189:CNPU7_7 port map (start_cn,clk,rst,V120C189,V499C189,V652C189,V678C189,V1065C189,V1341C189,V1437C189,C189V120,C189V499,C189V652,C189V678,C189V1065,C189V1341,C189V1437,end_cn189);
C190:CNPU7_7 port map (start_cn,clk,rst,V121C190,V500C190,V653C190,V679C190,V1066C190,V1342C190,V1438C190,C190V121,C190V500,C190V653,C190V679,C190V1066,C190V1342,C190V1438,end_cn190);
C191:CNPU7_7 port map (start_cn,clk,rst,V122C191,V501C191,V654C191,V680C191,V1067C191,V1343C191,V1439C191,C191V122,C191V501,C191V654,C191V680,C191V1067,C191V1343,C191V1439,end_cn191);
C192:CNPU7_7 port map (start_cn,clk,rst,V123C192,V502C192,V655C192,V681C192,V1068C192,V1344C192,V1440C192,C192V123,C192V502,C192V655,C192V681,C192V1068,C192V1344,C192V1440,end_cn192);
C193:CNPU7_7 port map (start_cn,clk,rst,V313C193,V407C193,V562C193,V706C193,V1057C193,V1345C193,V1441C193,C193V313,C193V407,C193V562,C193V706,C193V1057,C193V1345,C193V1441,end_cn193);
C194:CNPU7_7 port map (start_cn,clk,rst,V314C194,V408C194,V563C194,V707C194,V1058C194,V1346C194,V1442C194,C194V314,C194V408,C194V563,C194V707,C194V1058,C194V1346,C194V1442,end_cn194);
C195:CNPU7_7 port map (start_cn,clk,rst,V315C195,V409C195,V564C195,V708C195,V1059C195,V1347C195,V1443C195,C195V315,C195V409,C195V564,C195V708,C195V1059,C195V1347,C195V1443,end_cn195);
C196:CNPU7_7 port map (start_cn,clk,rst,V316C196,V410C196,V565C196,V709C196,V1060C196,V1348C196,V1444C196,C196V316,C196V410,C196V565,C196V709,C196V1060,C196V1348,C196V1444,end_cn196);
C197:CNPU7_7 port map (start_cn,clk,rst,V317C197,V411C197,V566C197,V710C197,V1061C197,V1349C197,V1445C197,C197V317,C197V411,C197V566,C197V710,C197V1061,C197V1349,C197V1445,end_cn197);
C198:CNPU7_7 port map (start_cn,clk,rst,V318C198,V412C198,V567C198,V711C198,V1062C198,V1350C198,V1446C198,C198V318,C198V412,C198V567,C198V711,C198V1062,C198V1350,C198V1446,end_cn198);
C199:CNPU7_7 port map (start_cn,clk,rst,V319C199,V413C199,V568C199,V712C199,V1063C199,V1351C199,V1447C199,C199V319,C199V413,C199V568,C199V712,C199V1063,C199V1351,C199V1447,end_cn199);
C200:CNPU7_7 port map (start_cn,clk,rst,V320C200,V414C200,V569C200,V713C200,V1064C200,V1352C200,V1448C200,C200V320,C200V414,C200V569,C200V713,C200V1064,C200V1352,C200V1448,end_cn200);
C201:CNPU7_7 port map (start_cn,clk,rst,V321C201,V415C201,V570C201,V714C201,V1065C201,V1353C201,V1449C201,C201V321,C201V415,C201V570,C201V714,C201V1065,C201V1353,C201V1449,end_cn201);
C202:CNPU7_7 port map (start_cn,clk,rst,V322C202,V416C202,V571C202,V715C202,V1066C202,V1354C202,V1450C202,C202V322,C202V416,C202V571,C202V715,C202V1066,C202V1354,C202V1450,end_cn202);
C203:CNPU7_7 port map (start_cn,clk,rst,V323C203,V417C203,V572C203,V716C203,V1067C203,V1355C203,V1451C203,C203V323,C203V417,C203V572,C203V716,C203V1067,C203V1355,C203V1451,end_cn203);
C204:CNPU7_7 port map (start_cn,clk,rst,V324C204,V418C204,V573C204,V717C204,V1068C204,V1356C204,V1452C204,C204V324,C204V418,C204V573,C204V717,C204V1068,C204V1356,C204V1452,end_cn204);
C205:CNPU7_7 port map (start_cn,clk,rst,V325C205,V419C205,V574C205,V718C205,V1069C205,V1357C205,V1453C205,C205V325,C205V419,C205V574,C205V718,C205V1069,C205V1357,C205V1453,end_cn205);
C206:CNPU7_7 port map (start_cn,clk,rst,V326C206,V420C206,V575C206,V719C206,V1070C206,V1358C206,V1454C206,C206V326,C206V420,C206V575,C206V719,C206V1070,C206V1358,C206V1454,end_cn206);
C207:CNPU7_7 port map (start_cn,clk,rst,V327C207,V421C207,V576C207,V720C207,V1071C207,V1359C207,V1455C207,C207V327,C207V421,C207V576,C207V720,C207V1071,C207V1359,C207V1455,end_cn207);
C208:CNPU7_7 port map (start_cn,clk,rst,V328C208,V422C208,V481C208,V721C208,V1072C208,V1360C208,V1456C208,C208V328,C208V422,C208V481,C208V721,C208V1072,C208V1360,C208V1456,end_cn208);
C209:CNPU7_7 port map (start_cn,clk,rst,V329C209,V423C209,V482C209,V722C209,V1073C209,V1361C209,V1457C209,C209V329,C209V423,C209V482,C209V722,C209V1073,C209V1361,C209V1457,end_cn209);
C210:CNPU7_7 port map (start_cn,clk,rst,V330C210,V424C210,V483C210,V723C210,V1074C210,V1362C210,V1458C210,C210V330,C210V424,C210V483,C210V723,C210V1074,C210V1362,C210V1458,end_cn210);
C211:CNPU7_7 port map (start_cn,clk,rst,V331C211,V425C211,V484C211,V724C211,V1075C211,V1363C211,V1459C211,C211V331,C211V425,C211V484,C211V724,C211V1075,C211V1363,C211V1459,end_cn211);
C212:CNPU7_7 port map (start_cn,clk,rst,V332C212,V426C212,V485C212,V725C212,V1076C212,V1364C212,V1460C212,C212V332,C212V426,C212V485,C212V725,C212V1076,C212V1364,C212V1460,end_cn212);
C213:CNPU7_7 port map (start_cn,clk,rst,V333C213,V427C213,V486C213,V726C213,V1077C213,V1365C213,V1461C213,C213V333,C213V427,C213V486,C213V726,C213V1077,C213V1365,C213V1461,end_cn213);
C214:CNPU7_7 port map (start_cn,clk,rst,V334C214,V428C214,V487C214,V727C214,V1078C214,V1366C214,V1462C214,C214V334,C214V428,C214V487,C214V727,C214V1078,C214V1366,C214V1462,end_cn214);
C215:CNPU7_7 port map (start_cn,clk,rst,V335C215,V429C215,V488C215,V728C215,V1079C215,V1367C215,V1463C215,C215V335,C215V429,C215V488,C215V728,C215V1079,C215V1367,C215V1463,end_cn215);
C216:CNPU7_7 port map (start_cn,clk,rst,V336C216,V430C216,V489C216,V729C216,V1080C216,V1368C216,V1464C216,C216V336,C216V430,C216V489,C216V729,C216V1080,C216V1368,C216V1464,end_cn216);
C217:CNPU7_7 port map (start_cn,clk,rst,V337C217,V431C217,V490C217,V730C217,V1081C217,V1369C217,V1465C217,C217V337,C217V431,C217V490,C217V730,C217V1081,C217V1369,C217V1465,end_cn217);
C218:CNPU7_7 port map (start_cn,clk,rst,V338C218,V432C218,V491C218,V731C218,V1082C218,V1370C218,V1466C218,C218V338,C218V432,C218V491,C218V731,C218V1082,C218V1370,C218V1466,end_cn218);
C219:CNPU7_7 port map (start_cn,clk,rst,V339C219,V433C219,V492C219,V732C219,V1083C219,V1371C219,V1467C219,C219V339,C219V433,C219V492,C219V732,C219V1083,C219V1371,C219V1467,end_cn219);
C220:CNPU7_7 port map (start_cn,clk,rst,V340C220,V434C220,V493C220,V733C220,V1084C220,V1372C220,V1468C220,C220V340,C220V434,C220V493,C220V733,C220V1084,C220V1372,C220V1468,end_cn220);
C221:CNPU7_7 port map (start_cn,clk,rst,V341C221,V435C221,V494C221,V734C221,V1085C221,V1373C221,V1469C221,C221V341,C221V435,C221V494,C221V734,C221V1085,C221V1373,C221V1469,end_cn221);
C222:CNPU7_7 port map (start_cn,clk,rst,V342C222,V436C222,V495C222,V735C222,V1086C222,V1374C222,V1470C222,C222V342,C222V436,C222V495,C222V735,C222V1086,C222V1374,C222V1470,end_cn222);
C223:CNPU7_7 port map (start_cn,clk,rst,V343C223,V437C223,V496C223,V736C223,V1087C223,V1375C223,V1471C223,C223V343,C223V437,C223V496,C223V736,C223V1087,C223V1375,C223V1471,end_cn223);
C224:CNPU7_7 port map (start_cn,clk,rst,V344C224,V438C224,V497C224,V737C224,V1088C224,V1376C224,V1472C224,C224V344,C224V438,C224V497,C224V737,C224V1088,C224V1376,C224V1472,end_cn224);
C225:CNPU7_7 port map (start_cn,clk,rst,V345C225,V439C225,V498C225,V738C225,V1089C225,V1377C225,V1473C225,C225V345,C225V439,C225V498,C225V738,C225V1089,C225V1377,C225V1473,end_cn225);
C226:CNPU7_7 port map (start_cn,clk,rst,V346C226,V440C226,V499C226,V739C226,V1090C226,V1378C226,V1474C226,C226V346,C226V440,C226V499,C226V739,C226V1090,C226V1378,C226V1474,end_cn226);
C227:CNPU7_7 port map (start_cn,clk,rst,V347C227,V441C227,V500C227,V740C227,V1091C227,V1379C227,V1475C227,C227V347,C227V441,C227V500,C227V740,C227V1091,C227V1379,C227V1475,end_cn227);
C228:CNPU7_7 port map (start_cn,clk,rst,V348C228,V442C228,V501C228,V741C228,V1092C228,V1380C228,V1476C228,C228V348,C228V442,C228V501,C228V741,C228V1092,C228V1380,C228V1476,end_cn228);
C229:CNPU7_7 port map (start_cn,clk,rst,V349C229,V443C229,V502C229,V742C229,V1093C229,V1381C229,V1477C229,C229V349,C229V443,C229V502,C229V742,C229V1093,C229V1381,C229V1477,end_cn229);
C230:CNPU7_7 port map (start_cn,clk,rst,V350C230,V444C230,V503C230,V743C230,V1094C230,V1382C230,V1478C230,C230V350,C230V444,C230V503,C230V743,C230V1094,C230V1382,C230V1478,end_cn230);
C231:CNPU7_7 port map (start_cn,clk,rst,V351C231,V445C231,V504C231,V744C231,V1095C231,V1383C231,V1479C231,C231V351,C231V445,C231V504,C231V744,C231V1095,C231V1383,C231V1479,end_cn231);
C232:CNPU7_7 port map (start_cn,clk,rst,V352C232,V446C232,V505C232,V745C232,V1096C232,V1384C232,V1480C232,C232V352,C232V446,C232V505,C232V745,C232V1096,C232V1384,C232V1480,end_cn232);
C233:CNPU7_7 port map (start_cn,clk,rst,V353C233,V447C233,V506C233,V746C233,V1097C233,V1385C233,V1481C233,C233V353,C233V447,C233V506,C233V746,C233V1097,C233V1385,C233V1481,end_cn233);
C234:CNPU7_7 port map (start_cn,clk,rst,V354C234,V448C234,V507C234,V747C234,V1098C234,V1386C234,V1482C234,C234V354,C234V448,C234V507,C234V747,C234V1098,C234V1386,C234V1482,end_cn234);
C235:CNPU7_7 port map (start_cn,clk,rst,V355C235,V449C235,V508C235,V748C235,V1099C235,V1387C235,V1483C235,C235V355,C235V449,C235V508,C235V748,C235V1099,C235V1387,C235V1483,end_cn235);
C236:CNPU7_7 port map (start_cn,clk,rst,V356C236,V450C236,V509C236,V749C236,V1100C236,V1388C236,V1484C236,C236V356,C236V450,C236V509,C236V749,C236V1100,C236V1388,C236V1484,end_cn236);
C237:CNPU7_7 port map (start_cn,clk,rst,V357C237,V451C237,V510C237,V750C237,V1101C237,V1389C237,V1485C237,C237V357,C237V451,C237V510,C237V750,C237V1101,C237V1389,C237V1485,end_cn237);
C238:CNPU7_7 port map (start_cn,clk,rst,V358C238,V452C238,V511C238,V751C238,V1102C238,V1390C238,V1486C238,C238V358,C238V452,C238V511,C238V751,C238V1102,C238V1390,C238V1486,end_cn238);
C239:CNPU7_7 port map (start_cn,clk,rst,V359C239,V453C239,V512C239,V752C239,V1103C239,V1391C239,V1487C239,C239V359,C239V453,C239V512,C239V752,C239V1103,C239V1391,C239V1487,end_cn239);
C240:CNPU7_7 port map (start_cn,clk,rst,V360C240,V454C240,V513C240,V753C240,V1104C240,V1392C240,V1488C240,C240V360,C240V454,C240V513,C240V753,C240V1104,C240V1392,C240V1488,end_cn240);
C241:CNPU7_7 port map (start_cn,clk,rst,V361C241,V455C241,V514C241,V754C241,V1105C241,V1393C241,V1489C241,C241V361,C241V455,C241V514,C241V754,C241V1105,C241V1393,C241V1489,end_cn241);
C242:CNPU7_7 port map (start_cn,clk,rst,V362C242,V456C242,V515C242,V755C242,V1106C242,V1394C242,V1490C242,C242V362,C242V456,C242V515,C242V755,C242V1106,C242V1394,C242V1490,end_cn242);
C243:CNPU7_7 port map (start_cn,clk,rst,V363C243,V457C243,V516C243,V756C243,V1107C243,V1395C243,V1491C243,C243V363,C243V457,C243V516,C243V756,C243V1107,C243V1395,C243V1491,end_cn243);
C244:CNPU7_7 port map (start_cn,clk,rst,V364C244,V458C244,V517C244,V757C244,V1108C244,V1396C244,V1492C244,C244V364,C244V458,C244V517,C244V757,C244V1108,C244V1396,C244V1492,end_cn244);
C245:CNPU7_7 port map (start_cn,clk,rst,V365C245,V459C245,V518C245,V758C245,V1109C245,V1397C245,V1493C245,C245V365,C245V459,C245V518,C245V758,C245V1109,C245V1397,C245V1493,end_cn245);
C246:CNPU7_7 port map (start_cn,clk,rst,V366C246,V460C246,V519C246,V759C246,V1110C246,V1398C246,V1494C246,C246V366,C246V460,C246V519,C246V759,C246V1110,C246V1398,C246V1494,end_cn246);
C247:CNPU7_7 port map (start_cn,clk,rst,V367C247,V461C247,V520C247,V760C247,V1111C247,V1399C247,V1495C247,C247V367,C247V461,C247V520,C247V760,C247V1111,C247V1399,C247V1495,end_cn247);
C248:CNPU7_7 port map (start_cn,clk,rst,V368C248,V462C248,V521C248,V761C248,V1112C248,V1400C248,V1496C248,C248V368,C248V462,C248V521,C248V761,C248V1112,C248V1400,C248V1496,end_cn248);
C249:CNPU7_7 port map (start_cn,clk,rst,V369C249,V463C249,V522C249,V762C249,V1113C249,V1401C249,V1497C249,C249V369,C249V463,C249V522,C249V762,C249V1113,C249V1401,C249V1497,end_cn249);
C250:CNPU7_7 port map (start_cn,clk,rst,V370C250,V464C250,V523C250,V763C250,V1114C250,V1402C250,V1498C250,C250V370,C250V464,C250V523,C250V763,C250V1114,C250V1402,C250V1498,end_cn250);
C251:CNPU7_7 port map (start_cn,clk,rst,V371C251,V465C251,V524C251,V764C251,V1115C251,V1403C251,V1499C251,C251V371,C251V465,C251V524,C251V764,C251V1115,C251V1403,C251V1499,end_cn251);
C252:CNPU7_7 port map (start_cn,clk,rst,V372C252,V466C252,V525C252,V765C252,V1116C252,V1404C252,V1500C252,C252V372,C252V466,C252V525,C252V765,C252V1116,C252V1404,C252V1500,end_cn252);
C253:CNPU7_7 port map (start_cn,clk,rst,V373C253,V467C253,V526C253,V766C253,V1117C253,V1405C253,V1501C253,C253V373,C253V467,C253V526,C253V766,C253V1117,C253V1405,C253V1501,end_cn253);
C254:CNPU7_7 port map (start_cn,clk,rst,V374C254,V468C254,V527C254,V767C254,V1118C254,V1406C254,V1502C254,C254V374,C254V468,C254V527,C254V767,C254V1118,C254V1406,C254V1502,end_cn254);
C255:CNPU7_7 port map (start_cn,clk,rst,V375C255,V469C255,V528C255,V768C255,V1119C255,V1407C255,V1503C255,C255V375,C255V469,C255V528,C255V768,C255V1119,C255V1407,C255V1503,end_cn255);
C256:CNPU7_7 port map (start_cn,clk,rst,V376C256,V470C256,V529C256,V673C256,V1120C256,V1408C256,V1504C256,C256V376,C256V470,C256V529,C256V673,C256V1120,C256V1408,C256V1504,end_cn256);
C257:CNPU7_7 port map (start_cn,clk,rst,V377C257,V471C257,V530C257,V674C257,V1121C257,V1409C257,V1505C257,C257V377,C257V471,C257V530,C257V674,C257V1121,C257V1409,C257V1505,end_cn257);
C258:CNPU7_7 port map (start_cn,clk,rst,V378C258,V472C258,V531C258,V675C258,V1122C258,V1410C258,V1506C258,C258V378,C258V472,C258V531,C258V675,C258V1122,C258V1410,C258V1506,end_cn258);
C259:CNPU7_7 port map (start_cn,clk,rst,V379C259,V473C259,V532C259,V676C259,V1123C259,V1411C259,V1507C259,C259V379,C259V473,C259V532,C259V676,C259V1123,C259V1411,C259V1507,end_cn259);
C260:CNPU7_7 port map (start_cn,clk,rst,V380C260,V474C260,V533C260,V677C260,V1124C260,V1412C260,V1508C260,C260V380,C260V474,C260V533,C260V677,C260V1124,C260V1412,C260V1508,end_cn260);
C261:CNPU7_7 port map (start_cn,clk,rst,V381C261,V475C261,V534C261,V678C261,V1125C261,V1413C261,V1509C261,C261V381,C261V475,C261V534,C261V678,C261V1125,C261V1413,C261V1509,end_cn261);
C262:CNPU7_7 port map (start_cn,clk,rst,V382C262,V476C262,V535C262,V679C262,V1126C262,V1414C262,V1510C262,C262V382,C262V476,C262V535,C262V679,C262V1126,C262V1414,C262V1510,end_cn262);
C263:CNPU7_7 port map (start_cn,clk,rst,V383C263,V477C263,V536C263,V680C263,V1127C263,V1415C263,V1511C263,C263V383,C263V477,C263V536,C263V680,C263V1127,C263V1415,C263V1511,end_cn263);
C264:CNPU7_7 port map (start_cn,clk,rst,V384C264,V478C264,V537C264,V681C264,V1128C264,V1416C264,V1512C264,C264V384,C264V478,C264V537,C264V681,C264V1128,C264V1416,C264V1512,end_cn264);
C265:CNPU7_7 port map (start_cn,clk,rst,V289C265,V479C265,V538C265,V682C265,V1129C265,V1417C265,V1513C265,C265V289,C265V479,C265V538,C265V682,C265V1129,C265V1417,C265V1513,end_cn265);
C266:CNPU7_7 port map (start_cn,clk,rst,V290C266,V480C266,V539C266,V683C266,V1130C266,V1418C266,V1514C266,C266V290,C266V480,C266V539,C266V683,C266V1130,C266V1418,C266V1514,end_cn266);
C267:CNPU7_7 port map (start_cn,clk,rst,V291C267,V385C267,V540C267,V684C267,V1131C267,V1419C267,V1515C267,C267V291,C267V385,C267V540,C267V684,C267V1131,C267V1419,C267V1515,end_cn267);
C268:CNPU7_7 port map (start_cn,clk,rst,V292C268,V386C268,V541C268,V685C268,V1132C268,V1420C268,V1516C268,C268V292,C268V386,C268V541,C268V685,C268V1132,C268V1420,C268V1516,end_cn268);
C269:CNPU7_7 port map (start_cn,clk,rst,V293C269,V387C269,V542C269,V686C269,V1133C269,V1421C269,V1517C269,C269V293,C269V387,C269V542,C269V686,C269V1133,C269V1421,C269V1517,end_cn269);
C270:CNPU7_7 port map (start_cn,clk,rst,V294C270,V388C270,V543C270,V687C270,V1134C270,V1422C270,V1518C270,C270V294,C270V388,C270V543,C270V687,C270V1134,C270V1422,C270V1518,end_cn270);
C271:CNPU7_7 port map (start_cn,clk,rst,V295C271,V389C271,V544C271,V688C271,V1135C271,V1423C271,V1519C271,C271V295,C271V389,C271V544,C271V688,C271V1135,C271V1423,C271V1519,end_cn271);
C272:CNPU7_7 port map (start_cn,clk,rst,V296C272,V390C272,V545C272,V689C272,V1136C272,V1424C272,V1520C272,C272V296,C272V390,C272V545,C272V689,C272V1136,C272V1424,C272V1520,end_cn272);
C273:CNPU7_7 port map (start_cn,clk,rst,V297C273,V391C273,V546C273,V690C273,V1137C273,V1425C273,V1521C273,C273V297,C273V391,C273V546,C273V690,C273V1137,C273V1425,C273V1521,end_cn273);
C274:CNPU7_7 port map (start_cn,clk,rst,V298C274,V392C274,V547C274,V691C274,V1138C274,V1426C274,V1522C274,C274V298,C274V392,C274V547,C274V691,C274V1138,C274V1426,C274V1522,end_cn274);
C275:CNPU7_7 port map (start_cn,clk,rst,V299C275,V393C275,V548C275,V692C275,V1139C275,V1427C275,V1523C275,C275V299,C275V393,C275V548,C275V692,C275V1139,C275V1427,C275V1523,end_cn275);
C276:CNPU7_7 port map (start_cn,clk,rst,V300C276,V394C276,V549C276,V693C276,V1140C276,V1428C276,V1524C276,C276V300,C276V394,C276V549,C276V693,C276V1140,C276V1428,C276V1524,end_cn276);
C277:CNPU7_7 port map (start_cn,clk,rst,V301C277,V395C277,V550C277,V694C277,V1141C277,V1429C277,V1525C277,C277V301,C277V395,C277V550,C277V694,C277V1141,C277V1429,C277V1525,end_cn277);
C278:CNPU7_7 port map (start_cn,clk,rst,V302C278,V396C278,V551C278,V695C278,V1142C278,V1430C278,V1526C278,C278V302,C278V396,C278V551,C278V695,C278V1142,C278V1430,C278V1526,end_cn278);
C279:CNPU7_7 port map (start_cn,clk,rst,V303C279,V397C279,V552C279,V696C279,V1143C279,V1431C279,V1527C279,C279V303,C279V397,C279V552,C279V696,C279V1143,C279V1431,C279V1527,end_cn279);
C280:CNPU7_7 port map (start_cn,clk,rst,V304C280,V398C280,V553C280,V697C280,V1144C280,V1432C280,V1528C280,C280V304,C280V398,C280V553,C280V697,C280V1144,C280V1432,C280V1528,end_cn280);
C281:CNPU7_7 port map (start_cn,clk,rst,V305C281,V399C281,V554C281,V698C281,V1145C281,V1433C281,V1529C281,C281V305,C281V399,C281V554,C281V698,C281V1145,C281V1433,C281V1529,end_cn281);
C282:CNPU7_7 port map (start_cn,clk,rst,V306C282,V400C282,V555C282,V699C282,V1146C282,V1434C282,V1530C282,C282V306,C282V400,C282V555,C282V699,C282V1146,C282V1434,C282V1530,end_cn282);
C283:CNPU7_7 port map (start_cn,clk,rst,V307C283,V401C283,V556C283,V700C283,V1147C283,V1435C283,V1531C283,C283V307,C283V401,C283V556,C283V700,C283V1147,C283V1435,C283V1531,end_cn283);
C284:CNPU7_7 port map (start_cn,clk,rst,V308C284,V402C284,V557C284,V701C284,V1148C284,V1436C284,V1532C284,C284V308,C284V402,C284V557,C284V701,C284V1148,C284V1436,C284V1532,end_cn284);
C285:CNPU7_7 port map (start_cn,clk,rst,V309C285,V403C285,V558C285,V702C285,V1149C285,V1437C285,V1533C285,C285V309,C285V403,C285V558,C285V702,C285V1149,C285V1437,C285V1533,end_cn285);
C286:CNPU7_7 port map (start_cn,clk,rst,V310C286,V404C286,V559C286,V703C286,V1150C286,V1438C286,V1534C286,C286V310,C286V404,C286V559,C286V703,C286V1150,C286V1438,C286V1534,end_cn286);
C287:CNPU7_7 port map (start_cn,clk,rst,V311C287,V405C287,V560C287,V704C287,V1151C287,V1439C287,V1535C287,C287V311,C287V405,C287V560,C287V704,C287V1151,C287V1439,C287V1535,end_cn287);
C288:CNPU7_7 port map (start_cn,clk,rst,V312C288,V406C288,V561C288,V705C288,V1152C288,V1440C288,V1536C288,C288V312,C288V406,C288V561,C288V705,C288V1152,C288V1440,C288V1536,end_cn288);
C289:CNPU6_6 port map (start_cn,clk,rst,V62C289,V240C289,V834C289,V890C289,V1441C289,V1537C289,C289V62,C289V240,C289V834,C289V890,C289V1441,C289V1537,end_cn289);
C290:CNPU6_6 port map (start_cn,clk,rst,V63C290,V241C290,V835C290,V891C290,V1442C290,V1538C290,C290V63,C290V241,C290V835,C290V891,C290V1442,C290V1538,end_cn290);
C291:CNPU6_6 port map (start_cn,clk,rst,V64C291,V242C291,V836C291,V892C291,V1443C291,V1539C291,C291V64,C291V242,C291V836,C291V892,C291V1443,C291V1539,end_cn291);
C292:CNPU6_6 port map (start_cn,clk,rst,V65C292,V243C292,V837C292,V893C292,V1444C292,V1540C292,C292V65,C292V243,C292V837,C292V893,C292V1444,C292V1540,end_cn292);
C293:CNPU6_6 port map (start_cn,clk,rst,V66C293,V244C293,V838C293,V894C293,V1445C293,V1541C293,C293V66,C293V244,C293V838,C293V894,C293V1445,C293V1541,end_cn293);
C294:CNPU6_6 port map (start_cn,clk,rst,V67C294,V245C294,V839C294,V895C294,V1446C294,V1542C294,C294V67,C294V245,C294V839,C294V895,C294V1446,C294V1542,end_cn294);
C295:CNPU6_6 port map (start_cn,clk,rst,V68C295,V246C295,V840C295,V896C295,V1447C295,V1543C295,C295V68,C295V246,C295V840,C295V896,C295V1447,C295V1543,end_cn295);
C296:CNPU6_6 port map (start_cn,clk,rst,V69C296,V247C296,V841C296,V897C296,V1448C296,V1544C296,C296V69,C296V247,C296V841,C296V897,C296V1448,C296V1544,end_cn296);
C297:CNPU6_6 port map (start_cn,clk,rst,V70C297,V248C297,V842C297,V898C297,V1449C297,V1545C297,C297V70,C297V248,C297V842,C297V898,C297V1449,C297V1545,end_cn297);
C298:CNPU6_6 port map (start_cn,clk,rst,V71C298,V249C298,V843C298,V899C298,V1450C298,V1546C298,C298V71,C298V249,C298V843,C298V899,C298V1450,C298V1546,end_cn298);
C299:CNPU6_6 port map (start_cn,clk,rst,V72C299,V250C299,V844C299,V900C299,V1451C299,V1547C299,C299V72,C299V250,C299V844,C299V900,C299V1451,C299V1547,end_cn299);
C300:CNPU6_6 port map (start_cn,clk,rst,V73C300,V251C300,V845C300,V901C300,V1452C300,V1548C300,C300V73,C300V251,C300V845,C300V901,C300V1452,C300V1548,end_cn300);
C301:CNPU6_6 port map (start_cn,clk,rst,V74C301,V252C301,V846C301,V902C301,V1453C301,V1549C301,C301V74,C301V252,C301V846,C301V902,C301V1453,C301V1549,end_cn301);
C302:CNPU6_6 port map (start_cn,clk,rst,V75C302,V253C302,V847C302,V903C302,V1454C302,V1550C302,C302V75,C302V253,C302V847,C302V903,C302V1454,C302V1550,end_cn302);
C303:CNPU6_6 port map (start_cn,clk,rst,V76C303,V254C303,V848C303,V904C303,V1455C303,V1551C303,C303V76,C303V254,C303V848,C303V904,C303V1455,C303V1551,end_cn303);
C304:CNPU6_6 port map (start_cn,clk,rst,V77C304,V255C304,V849C304,V905C304,V1456C304,V1552C304,C304V77,C304V255,C304V849,C304V905,C304V1456,C304V1552,end_cn304);
C305:CNPU6_6 port map (start_cn,clk,rst,V78C305,V256C305,V850C305,V906C305,V1457C305,V1553C305,C305V78,C305V256,C305V850,C305V906,C305V1457,C305V1553,end_cn305);
C306:CNPU6_6 port map (start_cn,clk,rst,V79C306,V257C306,V851C306,V907C306,V1458C306,V1554C306,C306V79,C306V257,C306V851,C306V907,C306V1458,C306V1554,end_cn306);
C307:CNPU6_6 port map (start_cn,clk,rst,V80C307,V258C307,V852C307,V908C307,V1459C307,V1555C307,C307V80,C307V258,C307V852,C307V908,C307V1459,C307V1555,end_cn307);
C308:CNPU6_6 port map (start_cn,clk,rst,V81C308,V259C308,V853C308,V909C308,V1460C308,V1556C308,C308V81,C308V259,C308V853,C308V909,C308V1460,C308V1556,end_cn308);
C309:CNPU6_6 port map (start_cn,clk,rst,V82C309,V260C309,V854C309,V910C309,V1461C309,V1557C309,C309V82,C309V260,C309V854,C309V910,C309V1461,C309V1557,end_cn309);
C310:CNPU6_6 port map (start_cn,clk,rst,V83C310,V261C310,V855C310,V911C310,V1462C310,V1558C310,C310V83,C310V261,C310V855,C310V911,C310V1462,C310V1558,end_cn310);
C311:CNPU6_6 port map (start_cn,clk,rst,V84C311,V262C311,V856C311,V912C311,V1463C311,V1559C311,C311V84,C311V262,C311V856,C311V912,C311V1463,C311V1559,end_cn311);
C312:CNPU6_6 port map (start_cn,clk,rst,V85C312,V263C312,V857C312,V913C312,V1464C312,V1560C312,C312V85,C312V263,C312V857,C312V913,C312V1464,C312V1560,end_cn312);
C313:CNPU6_6 port map (start_cn,clk,rst,V86C313,V264C313,V858C313,V914C313,V1465C313,V1561C313,C313V86,C313V264,C313V858,C313V914,C313V1465,C313V1561,end_cn313);
C314:CNPU6_6 port map (start_cn,clk,rst,V87C314,V265C314,V859C314,V915C314,V1466C314,V1562C314,C314V87,C314V265,C314V859,C314V915,C314V1466,C314V1562,end_cn314);
C315:CNPU6_6 port map (start_cn,clk,rst,V88C315,V266C315,V860C315,V916C315,V1467C315,V1563C315,C315V88,C315V266,C315V860,C315V916,C315V1467,C315V1563,end_cn315);
C316:CNPU6_6 port map (start_cn,clk,rst,V89C316,V267C316,V861C316,V917C316,V1468C316,V1564C316,C316V89,C316V267,C316V861,C316V917,C316V1468,C316V1564,end_cn316);
C317:CNPU6_6 port map (start_cn,clk,rst,V90C317,V268C317,V862C317,V918C317,V1469C317,V1565C317,C317V90,C317V268,C317V862,C317V918,C317V1469,C317V1565,end_cn317);
C318:CNPU6_6 port map (start_cn,clk,rst,V91C318,V269C318,V863C318,V919C318,V1470C318,V1566C318,C318V91,C318V269,C318V863,C318V919,C318V1470,C318V1566,end_cn318);
C319:CNPU6_6 port map (start_cn,clk,rst,V92C319,V270C319,V864C319,V920C319,V1471C319,V1567C319,C319V92,C319V270,C319V864,C319V920,C319V1471,C319V1567,end_cn319);
C320:CNPU6_6 port map (start_cn,clk,rst,V93C320,V271C320,V769C320,V921C320,V1472C320,V1568C320,C320V93,C320V271,C320V769,C320V921,C320V1472,C320V1568,end_cn320);
C321:CNPU6_6 port map (start_cn,clk,rst,V94C321,V272C321,V770C321,V922C321,V1473C321,V1569C321,C321V94,C321V272,C321V770,C321V922,C321V1473,C321V1569,end_cn321);
C322:CNPU6_6 port map (start_cn,clk,rst,V95C322,V273C322,V771C322,V923C322,V1474C322,V1570C322,C322V95,C322V273,C322V771,C322V923,C322V1474,C322V1570,end_cn322);
C323:CNPU6_6 port map (start_cn,clk,rst,V96C323,V274C323,V772C323,V924C323,V1475C323,V1571C323,C323V96,C323V274,C323V772,C323V924,C323V1475,C323V1571,end_cn323);
C324:CNPU6_6 port map (start_cn,clk,rst,V1C324,V275C324,V773C324,V925C324,V1476C324,V1572C324,C324V1,C324V275,C324V773,C324V925,C324V1476,C324V1572,end_cn324);
C325:CNPU6_6 port map (start_cn,clk,rst,V2C325,V276C325,V774C325,V926C325,V1477C325,V1573C325,C325V2,C325V276,C325V774,C325V926,C325V1477,C325V1573,end_cn325);
C326:CNPU6_6 port map (start_cn,clk,rst,V3C326,V277C326,V775C326,V927C326,V1478C326,V1574C326,C326V3,C326V277,C326V775,C326V927,C326V1478,C326V1574,end_cn326);
C327:CNPU6_6 port map (start_cn,clk,rst,V4C327,V278C327,V776C327,V928C327,V1479C327,V1575C327,C327V4,C327V278,C327V776,C327V928,C327V1479,C327V1575,end_cn327);
C328:CNPU6_6 port map (start_cn,clk,rst,V5C328,V279C328,V777C328,V929C328,V1480C328,V1576C328,C328V5,C328V279,C328V777,C328V929,C328V1480,C328V1576,end_cn328);
C329:CNPU6_6 port map (start_cn,clk,rst,V6C329,V280C329,V778C329,V930C329,V1481C329,V1577C329,C329V6,C329V280,C329V778,C329V930,C329V1481,C329V1577,end_cn329);
C330:CNPU6_6 port map (start_cn,clk,rst,V7C330,V281C330,V779C330,V931C330,V1482C330,V1578C330,C330V7,C330V281,C330V779,C330V931,C330V1482,C330V1578,end_cn330);
C331:CNPU6_6 port map (start_cn,clk,rst,V8C331,V282C331,V780C331,V932C331,V1483C331,V1579C331,C331V8,C331V282,C331V780,C331V932,C331V1483,C331V1579,end_cn331);
C332:CNPU6_6 port map (start_cn,clk,rst,V9C332,V283C332,V781C332,V933C332,V1484C332,V1580C332,C332V9,C332V283,C332V781,C332V933,C332V1484,C332V1580,end_cn332);
C333:CNPU6_6 port map (start_cn,clk,rst,V10C333,V284C333,V782C333,V934C333,V1485C333,V1581C333,C333V10,C333V284,C333V782,C333V934,C333V1485,C333V1581,end_cn333);
C334:CNPU6_6 port map (start_cn,clk,rst,V11C334,V285C334,V783C334,V935C334,V1486C334,V1582C334,C334V11,C334V285,C334V783,C334V935,C334V1486,C334V1582,end_cn334);
C335:CNPU6_6 port map (start_cn,clk,rst,V12C335,V286C335,V784C335,V936C335,V1487C335,V1583C335,C335V12,C335V286,C335V784,C335V936,C335V1487,C335V1583,end_cn335);
C336:CNPU6_6 port map (start_cn,clk,rst,V13C336,V287C336,V785C336,V937C336,V1488C336,V1584C336,C336V13,C336V287,C336V785,C336V937,C336V1488,C336V1584,end_cn336);
C337:CNPU6_6 port map (start_cn,clk,rst,V14C337,V288C337,V786C337,V938C337,V1489C337,V1585C337,C337V14,C337V288,C337V786,C337V938,C337V1489,C337V1585,end_cn337);
C338:CNPU6_6 port map (start_cn,clk,rst,V15C338,V193C338,V787C338,V939C338,V1490C338,V1586C338,C338V15,C338V193,C338V787,C338V939,C338V1490,C338V1586,end_cn338);
C339:CNPU6_6 port map (start_cn,clk,rst,V16C339,V194C339,V788C339,V940C339,V1491C339,V1587C339,C339V16,C339V194,C339V788,C339V940,C339V1491,C339V1587,end_cn339);
C340:CNPU6_6 port map (start_cn,clk,rst,V17C340,V195C340,V789C340,V941C340,V1492C340,V1588C340,C340V17,C340V195,C340V789,C340V941,C340V1492,C340V1588,end_cn340);
C341:CNPU6_6 port map (start_cn,clk,rst,V18C341,V196C341,V790C341,V942C341,V1493C341,V1589C341,C341V18,C341V196,C341V790,C341V942,C341V1493,C341V1589,end_cn341);
C342:CNPU6_6 port map (start_cn,clk,rst,V19C342,V197C342,V791C342,V943C342,V1494C342,V1590C342,C342V19,C342V197,C342V791,C342V943,C342V1494,C342V1590,end_cn342);
C343:CNPU6_6 port map (start_cn,clk,rst,V20C343,V198C343,V792C343,V944C343,V1495C343,V1591C343,C343V20,C343V198,C343V792,C343V944,C343V1495,C343V1591,end_cn343);
C344:CNPU6_6 port map (start_cn,clk,rst,V21C344,V199C344,V793C344,V945C344,V1496C344,V1592C344,C344V21,C344V199,C344V793,C344V945,C344V1496,C344V1592,end_cn344);
C345:CNPU6_6 port map (start_cn,clk,rst,V22C345,V200C345,V794C345,V946C345,V1497C345,V1593C345,C345V22,C345V200,C345V794,C345V946,C345V1497,C345V1593,end_cn345);
C346:CNPU6_6 port map (start_cn,clk,rst,V23C346,V201C346,V795C346,V947C346,V1498C346,V1594C346,C346V23,C346V201,C346V795,C346V947,C346V1498,C346V1594,end_cn346);
C347:CNPU6_6 port map (start_cn,clk,rst,V24C347,V202C347,V796C347,V948C347,V1499C347,V1595C347,C347V24,C347V202,C347V796,C347V948,C347V1499,C347V1595,end_cn347);
C348:CNPU6_6 port map (start_cn,clk,rst,V25C348,V203C348,V797C348,V949C348,V1500C348,V1596C348,C348V25,C348V203,C348V797,C348V949,C348V1500,C348V1596,end_cn348);
C349:CNPU6_6 port map (start_cn,clk,rst,V26C349,V204C349,V798C349,V950C349,V1501C349,V1597C349,C349V26,C349V204,C349V798,C349V950,C349V1501,C349V1597,end_cn349);
C350:CNPU6_6 port map (start_cn,clk,rst,V27C350,V205C350,V799C350,V951C350,V1502C350,V1598C350,C350V27,C350V205,C350V799,C350V951,C350V1502,C350V1598,end_cn350);
C351:CNPU6_6 port map (start_cn,clk,rst,V28C351,V206C351,V800C351,V952C351,V1503C351,V1599C351,C351V28,C351V206,C351V800,C351V952,C351V1503,C351V1599,end_cn351);
C352:CNPU6_6 port map (start_cn,clk,rst,V29C352,V207C352,V801C352,V953C352,V1504C352,V1600C352,C352V29,C352V207,C352V801,C352V953,C352V1504,C352V1600,end_cn352);
C353:CNPU6_6 port map (start_cn,clk,rst,V30C353,V208C353,V802C353,V954C353,V1505C353,V1601C353,C353V30,C353V208,C353V802,C353V954,C353V1505,C353V1601,end_cn353);
C354:CNPU6_6 port map (start_cn,clk,rst,V31C354,V209C354,V803C354,V955C354,V1506C354,V1602C354,C354V31,C354V209,C354V803,C354V955,C354V1506,C354V1602,end_cn354);
C355:CNPU6_6 port map (start_cn,clk,rst,V32C355,V210C355,V804C355,V956C355,V1507C355,V1603C355,C355V32,C355V210,C355V804,C355V956,C355V1507,C355V1603,end_cn355);
C356:CNPU6_6 port map (start_cn,clk,rst,V33C356,V211C356,V805C356,V957C356,V1508C356,V1604C356,C356V33,C356V211,C356V805,C356V957,C356V1508,C356V1604,end_cn356);
C357:CNPU6_6 port map (start_cn,clk,rst,V34C357,V212C357,V806C357,V958C357,V1509C357,V1605C357,C357V34,C357V212,C357V806,C357V958,C357V1509,C357V1605,end_cn357);
C358:CNPU6_6 port map (start_cn,clk,rst,V35C358,V213C358,V807C358,V959C358,V1510C358,V1606C358,C358V35,C358V213,C358V807,C358V959,C358V1510,C358V1606,end_cn358);
C359:CNPU6_6 port map (start_cn,clk,rst,V36C359,V214C359,V808C359,V960C359,V1511C359,V1607C359,C359V36,C359V214,C359V808,C359V960,C359V1511,C359V1607,end_cn359);
C360:CNPU6_6 port map (start_cn,clk,rst,V37C360,V215C360,V809C360,V865C360,V1512C360,V1608C360,C360V37,C360V215,C360V809,C360V865,C360V1512,C360V1608,end_cn360);
C361:CNPU6_6 port map (start_cn,clk,rst,V38C361,V216C361,V810C361,V866C361,V1513C361,V1609C361,C361V38,C361V216,C361V810,C361V866,C361V1513,C361V1609,end_cn361);
C362:CNPU6_6 port map (start_cn,clk,rst,V39C362,V217C362,V811C362,V867C362,V1514C362,V1610C362,C362V39,C362V217,C362V811,C362V867,C362V1514,C362V1610,end_cn362);
C363:CNPU6_6 port map (start_cn,clk,rst,V40C363,V218C363,V812C363,V868C363,V1515C363,V1611C363,C363V40,C363V218,C363V812,C363V868,C363V1515,C363V1611,end_cn363);
C364:CNPU6_6 port map (start_cn,clk,rst,V41C364,V219C364,V813C364,V869C364,V1516C364,V1612C364,C364V41,C364V219,C364V813,C364V869,C364V1516,C364V1612,end_cn364);
C365:CNPU6_6 port map (start_cn,clk,rst,V42C365,V220C365,V814C365,V870C365,V1517C365,V1613C365,C365V42,C365V220,C365V814,C365V870,C365V1517,C365V1613,end_cn365);
C366:CNPU6_6 port map (start_cn,clk,rst,V43C366,V221C366,V815C366,V871C366,V1518C366,V1614C366,C366V43,C366V221,C366V815,C366V871,C366V1518,C366V1614,end_cn366);
C367:CNPU6_6 port map (start_cn,clk,rst,V44C367,V222C367,V816C367,V872C367,V1519C367,V1615C367,C367V44,C367V222,C367V816,C367V872,C367V1519,C367V1615,end_cn367);
C368:CNPU6_6 port map (start_cn,clk,rst,V45C368,V223C368,V817C368,V873C368,V1520C368,V1616C368,C368V45,C368V223,C368V817,C368V873,C368V1520,C368V1616,end_cn368);
C369:CNPU6_6 port map (start_cn,clk,rst,V46C369,V224C369,V818C369,V874C369,V1521C369,V1617C369,C369V46,C369V224,C369V818,C369V874,C369V1521,C369V1617,end_cn369);
C370:CNPU6_6 port map (start_cn,clk,rst,V47C370,V225C370,V819C370,V875C370,V1522C370,V1618C370,C370V47,C370V225,C370V819,C370V875,C370V1522,C370V1618,end_cn370);
C371:CNPU6_6 port map (start_cn,clk,rst,V48C371,V226C371,V820C371,V876C371,V1523C371,V1619C371,C371V48,C371V226,C371V820,C371V876,C371V1523,C371V1619,end_cn371);
C372:CNPU6_6 port map (start_cn,clk,rst,V49C372,V227C372,V821C372,V877C372,V1524C372,V1620C372,C372V49,C372V227,C372V821,C372V877,C372V1524,C372V1620,end_cn372);
C373:CNPU6_6 port map (start_cn,clk,rst,V50C373,V228C373,V822C373,V878C373,V1525C373,V1621C373,C373V50,C373V228,C373V822,C373V878,C373V1525,C373V1621,end_cn373);
C374:CNPU6_6 port map (start_cn,clk,rst,V51C374,V229C374,V823C374,V879C374,V1526C374,V1622C374,C374V51,C374V229,C374V823,C374V879,C374V1526,C374V1622,end_cn374);
C375:CNPU6_6 port map (start_cn,clk,rst,V52C375,V230C375,V824C375,V880C375,V1527C375,V1623C375,C375V52,C375V230,C375V824,C375V880,C375V1527,C375V1623,end_cn375);
C376:CNPU6_6 port map (start_cn,clk,rst,V53C376,V231C376,V825C376,V881C376,V1528C376,V1624C376,C376V53,C376V231,C376V825,C376V881,C376V1528,C376V1624,end_cn376);
C377:CNPU6_6 port map (start_cn,clk,rst,V54C377,V232C377,V826C377,V882C377,V1529C377,V1625C377,C377V54,C377V232,C377V826,C377V882,C377V1529,C377V1625,end_cn377);
C378:CNPU6_6 port map (start_cn,clk,rst,V55C378,V233C378,V827C378,V883C378,V1530C378,V1626C378,C378V55,C378V233,C378V827,C378V883,C378V1530,C378V1626,end_cn378);
C379:CNPU6_6 port map (start_cn,clk,rst,V56C379,V234C379,V828C379,V884C379,V1531C379,V1627C379,C379V56,C379V234,C379V828,C379V884,C379V1531,C379V1627,end_cn379);
C380:CNPU6_6 port map (start_cn,clk,rst,V57C380,V235C380,V829C380,V885C380,V1532C380,V1628C380,C380V57,C380V235,C380V829,C380V885,C380V1532,C380V1628,end_cn380);
C381:CNPU6_6 port map (start_cn,clk,rst,V58C381,V236C381,V830C381,V886C381,V1533C381,V1629C381,C381V58,C381V236,C381V830,C381V886,C381V1533,C381V1629,end_cn381);
C382:CNPU6_6 port map (start_cn,clk,rst,V59C382,V237C382,V831C382,V887C382,V1534C382,V1630C382,C382V59,C382V237,C382V831,C382V887,C382V1534,C382V1630,end_cn382);
C383:CNPU6_6 port map (start_cn,clk,rst,V60C383,V238C383,V832C383,V888C383,V1535C383,V1631C383,C383V60,C383V238,C383V832,C383V888,C383V1535,C383V1631,end_cn383);
C384:CNPU6_6 port map (start_cn,clk,rst,V61C384,V239C384,V833C384,V889C384,V1536C384,V1632C384,C384V61,C384V239,C384V833,C384V889,C384V1536,C384V1632,end_cn384);
C385:CNPU6_6 port map (start_cn,clk,rst,V232C385,V661C385,V906C385,V1033C385,V1537C385,V1633C385,C385V232,C385V661,C385V906,C385V1033,C385V1537,C385V1633,end_cn385);
C386:CNPU6_6 port map (start_cn,clk,rst,V233C386,V662C386,V907C386,V1034C386,V1538C386,V1634C386,C386V233,C386V662,C386V907,C386V1034,C386V1538,C386V1634,end_cn386);
C387:CNPU6_6 port map (start_cn,clk,rst,V234C387,V663C387,V908C387,V1035C387,V1539C387,V1635C387,C387V234,C387V663,C387V908,C387V1035,C387V1539,C387V1635,end_cn387);
C388:CNPU6_6 port map (start_cn,clk,rst,V235C388,V664C388,V909C388,V1036C388,V1540C388,V1636C388,C388V235,C388V664,C388V909,C388V1036,C388V1540,C388V1636,end_cn388);
C389:CNPU6_6 port map (start_cn,clk,rst,V236C389,V665C389,V910C389,V1037C389,V1541C389,V1637C389,C389V236,C389V665,C389V910,C389V1037,C389V1541,C389V1637,end_cn389);
C390:CNPU6_6 port map (start_cn,clk,rst,V237C390,V666C390,V911C390,V1038C390,V1542C390,V1638C390,C390V237,C390V666,C390V911,C390V1038,C390V1542,C390V1638,end_cn390);
C391:CNPU6_6 port map (start_cn,clk,rst,V238C391,V667C391,V912C391,V1039C391,V1543C391,V1639C391,C391V238,C391V667,C391V912,C391V1039,C391V1543,C391V1639,end_cn391);
C392:CNPU6_6 port map (start_cn,clk,rst,V239C392,V668C392,V913C392,V1040C392,V1544C392,V1640C392,C392V239,C392V668,C392V913,C392V1040,C392V1544,C392V1640,end_cn392);
C393:CNPU6_6 port map (start_cn,clk,rst,V240C393,V669C393,V914C393,V1041C393,V1545C393,V1641C393,C393V240,C393V669,C393V914,C393V1041,C393V1545,C393V1641,end_cn393);
C394:CNPU6_6 port map (start_cn,clk,rst,V241C394,V670C394,V915C394,V1042C394,V1546C394,V1642C394,C394V241,C394V670,C394V915,C394V1042,C394V1546,C394V1642,end_cn394);
C395:CNPU6_6 port map (start_cn,clk,rst,V242C395,V671C395,V916C395,V1043C395,V1547C395,V1643C395,C395V242,C395V671,C395V916,C395V1043,C395V1547,C395V1643,end_cn395);
C396:CNPU6_6 port map (start_cn,clk,rst,V243C396,V672C396,V917C396,V1044C396,V1548C396,V1644C396,C396V243,C396V672,C396V917,C396V1044,C396V1548,C396V1644,end_cn396);
C397:CNPU6_6 port map (start_cn,clk,rst,V244C397,V577C397,V918C397,V1045C397,V1549C397,V1645C397,C397V244,C397V577,C397V918,C397V1045,C397V1549,C397V1645,end_cn397);
C398:CNPU6_6 port map (start_cn,clk,rst,V245C398,V578C398,V919C398,V1046C398,V1550C398,V1646C398,C398V245,C398V578,C398V919,C398V1046,C398V1550,C398V1646,end_cn398);
C399:CNPU6_6 port map (start_cn,clk,rst,V246C399,V579C399,V920C399,V1047C399,V1551C399,V1647C399,C399V246,C399V579,C399V920,C399V1047,C399V1551,C399V1647,end_cn399);
C400:CNPU6_6 port map (start_cn,clk,rst,V247C400,V580C400,V921C400,V1048C400,V1552C400,V1648C400,C400V247,C400V580,C400V921,C400V1048,C400V1552,C400V1648,end_cn400);
C401:CNPU6_6 port map (start_cn,clk,rst,V248C401,V581C401,V922C401,V1049C401,V1553C401,V1649C401,C401V248,C401V581,C401V922,C401V1049,C401V1553,C401V1649,end_cn401);
C402:CNPU6_6 port map (start_cn,clk,rst,V249C402,V582C402,V923C402,V1050C402,V1554C402,V1650C402,C402V249,C402V582,C402V923,C402V1050,C402V1554,C402V1650,end_cn402);
C403:CNPU6_6 port map (start_cn,clk,rst,V250C403,V583C403,V924C403,V1051C403,V1555C403,V1651C403,C403V250,C403V583,C403V924,C403V1051,C403V1555,C403V1651,end_cn403);
C404:CNPU6_6 port map (start_cn,clk,rst,V251C404,V584C404,V925C404,V1052C404,V1556C404,V1652C404,C404V251,C404V584,C404V925,C404V1052,C404V1556,C404V1652,end_cn404);
C405:CNPU6_6 port map (start_cn,clk,rst,V252C405,V585C405,V926C405,V1053C405,V1557C405,V1653C405,C405V252,C405V585,C405V926,C405V1053,C405V1557,C405V1653,end_cn405);
C406:CNPU6_6 port map (start_cn,clk,rst,V253C406,V586C406,V927C406,V1054C406,V1558C406,V1654C406,C406V253,C406V586,C406V927,C406V1054,C406V1558,C406V1654,end_cn406);
C407:CNPU6_6 port map (start_cn,clk,rst,V254C407,V587C407,V928C407,V1055C407,V1559C407,V1655C407,C407V254,C407V587,C407V928,C407V1055,C407V1559,C407V1655,end_cn407);
C408:CNPU6_6 port map (start_cn,clk,rst,V255C408,V588C408,V929C408,V1056C408,V1560C408,V1656C408,C408V255,C408V588,C408V929,C408V1056,C408V1560,C408V1656,end_cn408);
C409:CNPU6_6 port map (start_cn,clk,rst,V256C409,V589C409,V930C409,V961C409,V1561C409,V1657C409,C409V256,C409V589,C409V930,C409V961,C409V1561,C409V1657,end_cn409);
C410:CNPU6_6 port map (start_cn,clk,rst,V257C410,V590C410,V931C410,V962C410,V1562C410,V1658C410,C410V257,C410V590,C410V931,C410V962,C410V1562,C410V1658,end_cn410);
C411:CNPU6_6 port map (start_cn,clk,rst,V258C411,V591C411,V932C411,V963C411,V1563C411,V1659C411,C411V258,C411V591,C411V932,C411V963,C411V1563,C411V1659,end_cn411);
C412:CNPU6_6 port map (start_cn,clk,rst,V259C412,V592C412,V933C412,V964C412,V1564C412,V1660C412,C412V259,C412V592,C412V933,C412V964,C412V1564,C412V1660,end_cn412);
C413:CNPU6_6 port map (start_cn,clk,rst,V260C413,V593C413,V934C413,V965C413,V1565C413,V1661C413,C413V260,C413V593,C413V934,C413V965,C413V1565,C413V1661,end_cn413);
C414:CNPU6_6 port map (start_cn,clk,rst,V261C414,V594C414,V935C414,V966C414,V1566C414,V1662C414,C414V261,C414V594,C414V935,C414V966,C414V1566,C414V1662,end_cn414);
C415:CNPU6_6 port map (start_cn,clk,rst,V262C415,V595C415,V936C415,V967C415,V1567C415,V1663C415,C415V262,C415V595,C415V936,C415V967,C415V1567,C415V1663,end_cn415);
C416:CNPU6_6 port map (start_cn,clk,rst,V263C416,V596C416,V937C416,V968C416,V1568C416,V1664C416,C416V263,C416V596,C416V937,C416V968,C416V1568,C416V1664,end_cn416);
C417:CNPU6_6 port map (start_cn,clk,rst,V264C417,V597C417,V938C417,V969C417,V1569C417,V1665C417,C417V264,C417V597,C417V938,C417V969,C417V1569,C417V1665,end_cn417);
C418:CNPU6_6 port map (start_cn,clk,rst,V265C418,V598C418,V939C418,V970C418,V1570C418,V1666C418,C418V265,C418V598,C418V939,C418V970,C418V1570,C418V1666,end_cn418);
C419:CNPU6_6 port map (start_cn,clk,rst,V266C419,V599C419,V940C419,V971C419,V1571C419,V1667C419,C419V266,C419V599,C419V940,C419V971,C419V1571,C419V1667,end_cn419);
C420:CNPU6_6 port map (start_cn,clk,rst,V267C420,V600C420,V941C420,V972C420,V1572C420,V1668C420,C420V267,C420V600,C420V941,C420V972,C420V1572,C420V1668,end_cn420);
C421:CNPU6_6 port map (start_cn,clk,rst,V268C421,V601C421,V942C421,V973C421,V1573C421,V1669C421,C421V268,C421V601,C421V942,C421V973,C421V1573,C421V1669,end_cn421);
C422:CNPU6_6 port map (start_cn,clk,rst,V269C422,V602C422,V943C422,V974C422,V1574C422,V1670C422,C422V269,C422V602,C422V943,C422V974,C422V1574,C422V1670,end_cn422);
C423:CNPU6_6 port map (start_cn,clk,rst,V270C423,V603C423,V944C423,V975C423,V1575C423,V1671C423,C423V270,C423V603,C423V944,C423V975,C423V1575,C423V1671,end_cn423);
C424:CNPU6_6 port map (start_cn,clk,rst,V271C424,V604C424,V945C424,V976C424,V1576C424,V1672C424,C424V271,C424V604,C424V945,C424V976,C424V1576,C424V1672,end_cn424);
C425:CNPU6_6 port map (start_cn,clk,rst,V272C425,V605C425,V946C425,V977C425,V1577C425,V1673C425,C425V272,C425V605,C425V946,C425V977,C425V1577,C425V1673,end_cn425);
C426:CNPU6_6 port map (start_cn,clk,rst,V273C426,V606C426,V947C426,V978C426,V1578C426,V1674C426,C426V273,C426V606,C426V947,C426V978,C426V1578,C426V1674,end_cn426);
C427:CNPU6_6 port map (start_cn,clk,rst,V274C427,V607C427,V948C427,V979C427,V1579C427,V1675C427,C427V274,C427V607,C427V948,C427V979,C427V1579,C427V1675,end_cn427);
C428:CNPU6_6 port map (start_cn,clk,rst,V275C428,V608C428,V949C428,V980C428,V1580C428,V1676C428,C428V275,C428V608,C428V949,C428V980,C428V1580,C428V1676,end_cn428);
C429:CNPU6_6 port map (start_cn,clk,rst,V276C429,V609C429,V950C429,V981C429,V1581C429,V1677C429,C429V276,C429V609,C429V950,C429V981,C429V1581,C429V1677,end_cn429);
C430:CNPU6_6 port map (start_cn,clk,rst,V277C430,V610C430,V951C430,V982C430,V1582C430,V1678C430,C430V277,C430V610,C430V951,C430V982,C430V1582,C430V1678,end_cn430);
C431:CNPU6_6 port map (start_cn,clk,rst,V278C431,V611C431,V952C431,V983C431,V1583C431,V1679C431,C431V278,C431V611,C431V952,C431V983,C431V1583,C431V1679,end_cn431);
C432:CNPU6_6 port map (start_cn,clk,rst,V279C432,V612C432,V953C432,V984C432,V1584C432,V1680C432,C432V279,C432V612,C432V953,C432V984,C432V1584,C432V1680,end_cn432);
C433:CNPU6_6 port map (start_cn,clk,rst,V280C433,V613C433,V954C433,V985C433,V1585C433,V1681C433,C433V280,C433V613,C433V954,C433V985,C433V1585,C433V1681,end_cn433);
C434:CNPU6_6 port map (start_cn,clk,rst,V281C434,V614C434,V955C434,V986C434,V1586C434,V1682C434,C434V281,C434V614,C434V955,C434V986,C434V1586,C434V1682,end_cn434);
C435:CNPU6_6 port map (start_cn,clk,rst,V282C435,V615C435,V956C435,V987C435,V1587C435,V1683C435,C435V282,C435V615,C435V956,C435V987,C435V1587,C435V1683,end_cn435);
C436:CNPU6_6 port map (start_cn,clk,rst,V283C436,V616C436,V957C436,V988C436,V1588C436,V1684C436,C436V283,C436V616,C436V957,C436V988,C436V1588,C436V1684,end_cn436);
C437:CNPU6_6 port map (start_cn,clk,rst,V284C437,V617C437,V958C437,V989C437,V1589C437,V1685C437,C437V284,C437V617,C437V958,C437V989,C437V1589,C437V1685,end_cn437);
C438:CNPU6_6 port map (start_cn,clk,rst,V285C438,V618C438,V959C438,V990C438,V1590C438,V1686C438,C438V285,C438V618,C438V959,C438V990,C438V1590,C438V1686,end_cn438);
C439:CNPU6_6 port map (start_cn,clk,rst,V286C439,V619C439,V960C439,V991C439,V1591C439,V1687C439,C439V286,C439V619,C439V960,C439V991,C439V1591,C439V1687,end_cn439);
C440:CNPU6_6 port map (start_cn,clk,rst,V287C440,V620C440,V865C440,V992C440,V1592C440,V1688C440,C440V287,C440V620,C440V865,C440V992,C440V1592,C440V1688,end_cn440);
C441:CNPU6_6 port map (start_cn,clk,rst,V288C441,V621C441,V866C441,V993C441,V1593C441,V1689C441,C441V288,C441V621,C441V866,C441V993,C441V1593,C441V1689,end_cn441);
C442:CNPU6_6 port map (start_cn,clk,rst,V193C442,V622C442,V867C442,V994C442,V1594C442,V1690C442,C442V193,C442V622,C442V867,C442V994,C442V1594,C442V1690,end_cn442);
C443:CNPU6_6 port map (start_cn,clk,rst,V194C443,V623C443,V868C443,V995C443,V1595C443,V1691C443,C443V194,C443V623,C443V868,C443V995,C443V1595,C443V1691,end_cn443);
C444:CNPU6_6 port map (start_cn,clk,rst,V195C444,V624C444,V869C444,V996C444,V1596C444,V1692C444,C444V195,C444V624,C444V869,C444V996,C444V1596,C444V1692,end_cn444);
C445:CNPU6_6 port map (start_cn,clk,rst,V196C445,V625C445,V870C445,V997C445,V1597C445,V1693C445,C445V196,C445V625,C445V870,C445V997,C445V1597,C445V1693,end_cn445);
C446:CNPU6_6 port map (start_cn,clk,rst,V197C446,V626C446,V871C446,V998C446,V1598C446,V1694C446,C446V197,C446V626,C446V871,C446V998,C446V1598,C446V1694,end_cn446);
C447:CNPU6_6 port map (start_cn,clk,rst,V198C447,V627C447,V872C447,V999C447,V1599C447,V1695C447,C447V198,C447V627,C447V872,C447V999,C447V1599,C447V1695,end_cn447);
C448:CNPU6_6 port map (start_cn,clk,rst,V199C448,V628C448,V873C448,V1000C448,V1600C448,V1696C448,C448V199,C448V628,C448V873,C448V1000,C448V1600,C448V1696,end_cn448);
C449:CNPU6_6 port map (start_cn,clk,rst,V200C449,V629C449,V874C449,V1001C449,V1601C449,V1697C449,C449V200,C449V629,C449V874,C449V1001,C449V1601,C449V1697,end_cn449);
C450:CNPU6_6 port map (start_cn,clk,rst,V201C450,V630C450,V875C450,V1002C450,V1602C450,V1698C450,C450V201,C450V630,C450V875,C450V1002,C450V1602,C450V1698,end_cn450);
C451:CNPU6_6 port map (start_cn,clk,rst,V202C451,V631C451,V876C451,V1003C451,V1603C451,V1699C451,C451V202,C451V631,C451V876,C451V1003,C451V1603,C451V1699,end_cn451);
C452:CNPU6_6 port map (start_cn,clk,rst,V203C452,V632C452,V877C452,V1004C452,V1604C452,V1700C452,C452V203,C452V632,C452V877,C452V1004,C452V1604,C452V1700,end_cn452);
C453:CNPU6_6 port map (start_cn,clk,rst,V204C453,V633C453,V878C453,V1005C453,V1605C453,V1701C453,C453V204,C453V633,C453V878,C453V1005,C453V1605,C453V1701,end_cn453);
C454:CNPU6_6 port map (start_cn,clk,rst,V205C454,V634C454,V879C454,V1006C454,V1606C454,V1702C454,C454V205,C454V634,C454V879,C454V1006,C454V1606,C454V1702,end_cn454);
C455:CNPU6_6 port map (start_cn,clk,rst,V206C455,V635C455,V880C455,V1007C455,V1607C455,V1703C455,C455V206,C455V635,C455V880,C455V1007,C455V1607,C455V1703,end_cn455);
C456:CNPU6_6 port map (start_cn,clk,rst,V207C456,V636C456,V881C456,V1008C456,V1608C456,V1704C456,C456V207,C456V636,C456V881,C456V1008,C456V1608,C456V1704,end_cn456);
C457:CNPU6_6 port map (start_cn,clk,rst,V208C457,V637C457,V882C457,V1009C457,V1609C457,V1705C457,C457V208,C457V637,C457V882,C457V1009,C457V1609,C457V1705,end_cn457);
C458:CNPU6_6 port map (start_cn,clk,rst,V209C458,V638C458,V883C458,V1010C458,V1610C458,V1706C458,C458V209,C458V638,C458V883,C458V1010,C458V1610,C458V1706,end_cn458);
C459:CNPU6_6 port map (start_cn,clk,rst,V210C459,V639C459,V884C459,V1011C459,V1611C459,V1707C459,C459V210,C459V639,C459V884,C459V1011,C459V1611,C459V1707,end_cn459);
C460:CNPU6_6 port map (start_cn,clk,rst,V211C460,V640C460,V885C460,V1012C460,V1612C460,V1708C460,C460V211,C460V640,C460V885,C460V1012,C460V1612,C460V1708,end_cn460);
C461:CNPU6_6 port map (start_cn,clk,rst,V212C461,V641C461,V886C461,V1013C461,V1613C461,V1709C461,C461V212,C461V641,C461V886,C461V1013,C461V1613,C461V1709,end_cn461);
C462:CNPU6_6 port map (start_cn,clk,rst,V213C462,V642C462,V887C462,V1014C462,V1614C462,V1710C462,C462V213,C462V642,C462V887,C462V1014,C462V1614,C462V1710,end_cn462);
C463:CNPU6_6 port map (start_cn,clk,rst,V214C463,V643C463,V888C463,V1015C463,V1615C463,V1711C463,C463V214,C463V643,C463V888,C463V1015,C463V1615,C463V1711,end_cn463);
C464:CNPU6_6 port map (start_cn,clk,rst,V215C464,V644C464,V889C464,V1016C464,V1616C464,V1712C464,C464V215,C464V644,C464V889,C464V1016,C464V1616,C464V1712,end_cn464);
C465:CNPU6_6 port map (start_cn,clk,rst,V216C465,V645C465,V890C465,V1017C465,V1617C465,V1713C465,C465V216,C465V645,C465V890,C465V1017,C465V1617,C465V1713,end_cn465);
C466:CNPU6_6 port map (start_cn,clk,rst,V217C466,V646C466,V891C466,V1018C466,V1618C466,V1714C466,C466V217,C466V646,C466V891,C466V1018,C466V1618,C466V1714,end_cn466);
C467:CNPU6_6 port map (start_cn,clk,rst,V218C467,V647C467,V892C467,V1019C467,V1619C467,V1715C467,C467V218,C467V647,C467V892,C467V1019,C467V1619,C467V1715,end_cn467);
C468:CNPU6_6 port map (start_cn,clk,rst,V219C468,V648C468,V893C468,V1020C468,V1620C468,V1716C468,C468V219,C468V648,C468V893,C468V1020,C468V1620,C468V1716,end_cn468);
C469:CNPU6_6 port map (start_cn,clk,rst,V220C469,V649C469,V894C469,V1021C469,V1621C469,V1717C469,C469V220,C469V649,C469V894,C469V1021,C469V1621,C469V1717,end_cn469);
C470:CNPU6_6 port map (start_cn,clk,rst,V221C470,V650C470,V895C470,V1022C470,V1622C470,V1718C470,C470V221,C470V650,C470V895,C470V1022,C470V1622,C470V1718,end_cn470);
C471:CNPU6_6 port map (start_cn,clk,rst,V222C471,V651C471,V896C471,V1023C471,V1623C471,V1719C471,C471V222,C471V651,C471V896,C471V1023,C471V1623,C471V1719,end_cn471);
C472:CNPU6_6 port map (start_cn,clk,rst,V223C472,V652C472,V897C472,V1024C472,V1624C472,V1720C472,C472V223,C472V652,C472V897,C472V1024,C472V1624,C472V1720,end_cn472);
C473:CNPU6_6 port map (start_cn,clk,rst,V224C473,V653C473,V898C473,V1025C473,V1625C473,V1721C473,C473V224,C473V653,C473V898,C473V1025,C473V1625,C473V1721,end_cn473);
C474:CNPU6_6 port map (start_cn,clk,rst,V225C474,V654C474,V899C474,V1026C474,V1626C474,V1722C474,C474V225,C474V654,C474V899,C474V1026,C474V1626,C474V1722,end_cn474);
C475:CNPU6_6 port map (start_cn,clk,rst,V226C475,V655C475,V900C475,V1027C475,V1627C475,V1723C475,C475V226,C475V655,C475V900,C475V1027,C475V1627,C475V1723,end_cn475);
C476:CNPU6_6 port map (start_cn,clk,rst,V227C476,V656C476,V901C476,V1028C476,V1628C476,V1724C476,C476V227,C476V656,C476V901,C476V1028,C476V1628,C476V1724,end_cn476);
C477:CNPU6_6 port map (start_cn,clk,rst,V228C477,V657C477,V902C477,V1029C477,V1629C477,V1725C477,C477V228,C477V657,C477V902,C477V1029,C477V1629,C477V1725,end_cn477);
C478:CNPU6_6 port map (start_cn,clk,rst,V229C478,V658C478,V903C478,V1030C478,V1630C478,V1726C478,C478V229,C478V658,C478V903,C478V1030,C478V1630,C478V1726,end_cn478);
C479:CNPU6_6 port map (start_cn,clk,rst,V230C479,V659C479,V904C479,V1031C479,V1631C479,V1727C479,C479V230,C479V659,C479V904,C479V1031,C479V1631,C479V1727,end_cn479);
C480:CNPU6_6 port map (start_cn,clk,rst,V231C480,V660C480,V905C480,V1032C480,V1632C480,V1728C480,C480V231,C480V660,C480V905,C480V1032,C480V1632,C480V1728,end_cn480);
C481:CNPU7_7 port map (start_cn,clk,rst,V431C481,V521C481,V755C481,V1136C481,V1153C481,V1633C481,V1729C481,C481V431,C481V521,C481V755,C481V1136,C481V1153,C481V1633,C481V1729,end_cn481);
C482:CNPU7_7 port map (start_cn,clk,rst,V432C482,V522C482,V756C482,V1137C482,V1154C482,V1634C482,V1730C482,C482V432,C482V522,C482V756,C482V1137,C482V1154,C482V1634,C482V1730,end_cn482);
C483:CNPU7_7 port map (start_cn,clk,rst,V433C483,V523C483,V757C483,V1138C483,V1155C483,V1635C483,V1731C483,C483V433,C483V523,C483V757,C483V1138,C483V1155,C483V1635,C483V1731,end_cn483);
C484:CNPU7_7 port map (start_cn,clk,rst,V434C484,V524C484,V758C484,V1139C484,V1156C484,V1636C484,V1732C484,C484V434,C484V524,C484V758,C484V1139,C484V1156,C484V1636,C484V1732,end_cn484);
C485:CNPU7_7 port map (start_cn,clk,rst,V435C485,V525C485,V759C485,V1140C485,V1157C485,V1637C485,V1733C485,C485V435,C485V525,C485V759,C485V1140,C485V1157,C485V1637,C485V1733,end_cn485);
C486:CNPU7_7 port map (start_cn,clk,rst,V436C486,V526C486,V760C486,V1141C486,V1158C486,V1638C486,V1734C486,C486V436,C486V526,C486V760,C486V1141,C486V1158,C486V1638,C486V1734,end_cn486);
C487:CNPU7_7 port map (start_cn,clk,rst,V437C487,V527C487,V761C487,V1142C487,V1159C487,V1639C487,V1735C487,C487V437,C487V527,C487V761,C487V1142,C487V1159,C487V1639,C487V1735,end_cn487);
C488:CNPU7_7 port map (start_cn,clk,rst,V438C488,V528C488,V762C488,V1143C488,V1160C488,V1640C488,V1736C488,C488V438,C488V528,C488V762,C488V1143,C488V1160,C488V1640,C488V1736,end_cn488);
C489:CNPU7_7 port map (start_cn,clk,rst,V439C489,V529C489,V763C489,V1144C489,V1161C489,V1641C489,V1737C489,C489V439,C489V529,C489V763,C489V1144,C489V1161,C489V1641,C489V1737,end_cn489);
C490:CNPU7_7 port map (start_cn,clk,rst,V440C490,V530C490,V764C490,V1145C490,V1162C490,V1642C490,V1738C490,C490V440,C490V530,C490V764,C490V1145,C490V1162,C490V1642,C490V1738,end_cn490);
C491:CNPU7_7 port map (start_cn,clk,rst,V441C491,V531C491,V765C491,V1146C491,V1163C491,V1643C491,V1739C491,C491V441,C491V531,C491V765,C491V1146,C491V1163,C491V1643,C491V1739,end_cn491);
C492:CNPU7_7 port map (start_cn,clk,rst,V442C492,V532C492,V766C492,V1147C492,V1164C492,V1644C492,V1740C492,C492V442,C492V532,C492V766,C492V1147,C492V1164,C492V1644,C492V1740,end_cn492);
C493:CNPU7_7 port map (start_cn,clk,rst,V443C493,V533C493,V767C493,V1148C493,V1165C493,V1645C493,V1741C493,C493V443,C493V533,C493V767,C493V1148,C493V1165,C493V1645,C493V1741,end_cn493);
C494:CNPU7_7 port map (start_cn,clk,rst,V444C494,V534C494,V768C494,V1149C494,V1166C494,V1646C494,V1742C494,C494V444,C494V534,C494V768,C494V1149,C494V1166,C494V1646,C494V1742,end_cn494);
C495:CNPU7_7 port map (start_cn,clk,rst,V445C495,V535C495,V673C495,V1150C495,V1167C495,V1647C495,V1743C495,C495V445,C495V535,C495V673,C495V1150,C495V1167,C495V1647,C495V1743,end_cn495);
C496:CNPU7_7 port map (start_cn,clk,rst,V446C496,V536C496,V674C496,V1151C496,V1168C496,V1648C496,V1744C496,C496V446,C496V536,C496V674,C496V1151,C496V1168,C496V1648,C496V1744,end_cn496);
C497:CNPU7_7 port map (start_cn,clk,rst,V447C497,V537C497,V675C497,V1152C497,V1169C497,V1649C497,V1745C497,C497V447,C497V537,C497V675,C497V1152,C497V1169,C497V1649,C497V1745,end_cn497);
C498:CNPU7_7 port map (start_cn,clk,rst,V448C498,V538C498,V676C498,V1057C498,V1170C498,V1650C498,V1746C498,C498V448,C498V538,C498V676,C498V1057,C498V1170,C498V1650,C498V1746,end_cn498);
C499:CNPU7_7 port map (start_cn,clk,rst,V449C499,V539C499,V677C499,V1058C499,V1171C499,V1651C499,V1747C499,C499V449,C499V539,C499V677,C499V1058,C499V1171,C499V1651,C499V1747,end_cn499);
C500:CNPU7_7 port map (start_cn,clk,rst,V450C500,V540C500,V678C500,V1059C500,V1172C500,V1652C500,V1748C500,C500V450,C500V540,C500V678,C500V1059,C500V1172,C500V1652,C500V1748,end_cn500);
C501:CNPU7_7 port map (start_cn,clk,rst,V451C501,V541C501,V679C501,V1060C501,V1173C501,V1653C501,V1749C501,C501V451,C501V541,C501V679,C501V1060,C501V1173,C501V1653,C501V1749,end_cn501);
C502:CNPU7_7 port map (start_cn,clk,rst,V452C502,V542C502,V680C502,V1061C502,V1174C502,V1654C502,V1750C502,C502V452,C502V542,C502V680,C502V1061,C502V1174,C502V1654,C502V1750,end_cn502);
C503:CNPU7_7 port map (start_cn,clk,rst,V453C503,V543C503,V681C503,V1062C503,V1175C503,V1655C503,V1751C503,C503V453,C503V543,C503V681,C503V1062,C503V1175,C503V1655,C503V1751,end_cn503);
C504:CNPU7_7 port map (start_cn,clk,rst,V454C504,V544C504,V682C504,V1063C504,V1176C504,V1656C504,V1752C504,C504V454,C504V544,C504V682,C504V1063,C504V1176,C504V1656,C504V1752,end_cn504);
C505:CNPU7_7 port map (start_cn,clk,rst,V455C505,V545C505,V683C505,V1064C505,V1177C505,V1657C505,V1753C505,C505V455,C505V545,C505V683,C505V1064,C505V1177,C505V1657,C505V1753,end_cn505);
C506:CNPU7_7 port map (start_cn,clk,rst,V456C506,V546C506,V684C506,V1065C506,V1178C506,V1658C506,V1754C506,C506V456,C506V546,C506V684,C506V1065,C506V1178,C506V1658,C506V1754,end_cn506);
C507:CNPU7_7 port map (start_cn,clk,rst,V457C507,V547C507,V685C507,V1066C507,V1179C507,V1659C507,V1755C507,C507V457,C507V547,C507V685,C507V1066,C507V1179,C507V1659,C507V1755,end_cn507);
C508:CNPU7_7 port map (start_cn,clk,rst,V458C508,V548C508,V686C508,V1067C508,V1180C508,V1660C508,V1756C508,C508V458,C508V548,C508V686,C508V1067,C508V1180,C508V1660,C508V1756,end_cn508);
C509:CNPU7_7 port map (start_cn,clk,rst,V459C509,V549C509,V687C509,V1068C509,V1181C509,V1661C509,V1757C509,C509V459,C509V549,C509V687,C509V1068,C509V1181,C509V1661,C509V1757,end_cn509);
C510:CNPU7_7 port map (start_cn,clk,rst,V460C510,V550C510,V688C510,V1069C510,V1182C510,V1662C510,V1758C510,C510V460,C510V550,C510V688,C510V1069,C510V1182,C510V1662,C510V1758,end_cn510);
C511:CNPU7_7 port map (start_cn,clk,rst,V461C511,V551C511,V689C511,V1070C511,V1183C511,V1663C511,V1759C511,C511V461,C511V551,C511V689,C511V1070,C511V1183,C511V1663,C511V1759,end_cn511);
C512:CNPU7_7 port map (start_cn,clk,rst,V462C512,V552C512,V690C512,V1071C512,V1184C512,V1664C512,V1760C512,C512V462,C512V552,C512V690,C512V1071,C512V1184,C512V1664,C512V1760,end_cn512);
C513:CNPU7_7 port map (start_cn,clk,rst,V463C513,V553C513,V691C513,V1072C513,V1185C513,V1665C513,V1761C513,C513V463,C513V553,C513V691,C513V1072,C513V1185,C513V1665,C513V1761,end_cn513);
C514:CNPU7_7 port map (start_cn,clk,rst,V464C514,V554C514,V692C514,V1073C514,V1186C514,V1666C514,V1762C514,C514V464,C514V554,C514V692,C514V1073,C514V1186,C514V1666,C514V1762,end_cn514);
C515:CNPU7_7 port map (start_cn,clk,rst,V465C515,V555C515,V693C515,V1074C515,V1187C515,V1667C515,V1763C515,C515V465,C515V555,C515V693,C515V1074,C515V1187,C515V1667,C515V1763,end_cn515);
C516:CNPU7_7 port map (start_cn,clk,rst,V466C516,V556C516,V694C516,V1075C516,V1188C516,V1668C516,V1764C516,C516V466,C516V556,C516V694,C516V1075,C516V1188,C516V1668,C516V1764,end_cn516);
C517:CNPU7_7 port map (start_cn,clk,rst,V467C517,V557C517,V695C517,V1076C517,V1189C517,V1669C517,V1765C517,C517V467,C517V557,C517V695,C517V1076,C517V1189,C517V1669,C517V1765,end_cn517);
C518:CNPU7_7 port map (start_cn,clk,rst,V468C518,V558C518,V696C518,V1077C518,V1190C518,V1670C518,V1766C518,C518V468,C518V558,C518V696,C518V1077,C518V1190,C518V1670,C518V1766,end_cn518);
C519:CNPU7_7 port map (start_cn,clk,rst,V469C519,V559C519,V697C519,V1078C519,V1191C519,V1671C519,V1767C519,C519V469,C519V559,C519V697,C519V1078,C519V1191,C519V1671,C519V1767,end_cn519);
C520:CNPU7_7 port map (start_cn,clk,rst,V470C520,V560C520,V698C520,V1079C520,V1192C520,V1672C520,V1768C520,C520V470,C520V560,C520V698,C520V1079,C520V1192,C520V1672,C520V1768,end_cn520);
C521:CNPU7_7 port map (start_cn,clk,rst,V471C521,V561C521,V699C521,V1080C521,V1193C521,V1673C521,V1769C521,C521V471,C521V561,C521V699,C521V1080,C521V1193,C521V1673,C521V1769,end_cn521);
C522:CNPU7_7 port map (start_cn,clk,rst,V472C522,V562C522,V700C522,V1081C522,V1194C522,V1674C522,V1770C522,C522V472,C522V562,C522V700,C522V1081,C522V1194,C522V1674,C522V1770,end_cn522);
C523:CNPU7_7 port map (start_cn,clk,rst,V473C523,V563C523,V701C523,V1082C523,V1195C523,V1675C523,V1771C523,C523V473,C523V563,C523V701,C523V1082,C523V1195,C523V1675,C523V1771,end_cn523);
C524:CNPU7_7 port map (start_cn,clk,rst,V474C524,V564C524,V702C524,V1083C524,V1196C524,V1676C524,V1772C524,C524V474,C524V564,C524V702,C524V1083,C524V1196,C524V1676,C524V1772,end_cn524);
C525:CNPU7_7 port map (start_cn,clk,rst,V475C525,V565C525,V703C525,V1084C525,V1197C525,V1677C525,V1773C525,C525V475,C525V565,C525V703,C525V1084,C525V1197,C525V1677,C525V1773,end_cn525);
C526:CNPU7_7 port map (start_cn,clk,rst,V476C526,V566C526,V704C526,V1085C526,V1198C526,V1678C526,V1774C526,C526V476,C526V566,C526V704,C526V1085,C526V1198,C526V1678,C526V1774,end_cn526);
C527:CNPU7_7 port map (start_cn,clk,rst,V477C527,V567C527,V705C527,V1086C527,V1199C527,V1679C527,V1775C527,C527V477,C527V567,C527V705,C527V1086,C527V1199,C527V1679,C527V1775,end_cn527);
C528:CNPU7_7 port map (start_cn,clk,rst,V478C528,V568C528,V706C528,V1087C528,V1200C528,V1680C528,V1776C528,C528V478,C528V568,C528V706,C528V1087,C528V1200,C528V1680,C528V1776,end_cn528);
C529:CNPU7_7 port map (start_cn,clk,rst,V479C529,V569C529,V707C529,V1088C529,V1201C529,V1681C529,V1777C529,C529V479,C529V569,C529V707,C529V1088,C529V1201,C529V1681,C529V1777,end_cn529);
C530:CNPU7_7 port map (start_cn,clk,rst,V480C530,V570C530,V708C530,V1089C530,V1202C530,V1682C530,V1778C530,C530V480,C530V570,C530V708,C530V1089,C530V1202,C530V1682,C530V1778,end_cn530);
C531:CNPU7_7 port map (start_cn,clk,rst,V385C531,V571C531,V709C531,V1090C531,V1203C531,V1683C531,V1779C531,C531V385,C531V571,C531V709,C531V1090,C531V1203,C531V1683,C531V1779,end_cn531);
C532:CNPU7_7 port map (start_cn,clk,rst,V386C532,V572C532,V710C532,V1091C532,V1204C532,V1684C532,V1780C532,C532V386,C532V572,C532V710,C532V1091,C532V1204,C532V1684,C532V1780,end_cn532);
C533:CNPU7_7 port map (start_cn,clk,rst,V387C533,V573C533,V711C533,V1092C533,V1205C533,V1685C533,V1781C533,C533V387,C533V573,C533V711,C533V1092,C533V1205,C533V1685,C533V1781,end_cn533);
C534:CNPU7_7 port map (start_cn,clk,rst,V388C534,V574C534,V712C534,V1093C534,V1206C534,V1686C534,V1782C534,C534V388,C534V574,C534V712,C534V1093,C534V1206,C534V1686,C534V1782,end_cn534);
C535:CNPU7_7 port map (start_cn,clk,rst,V389C535,V575C535,V713C535,V1094C535,V1207C535,V1687C535,V1783C535,C535V389,C535V575,C535V713,C535V1094,C535V1207,C535V1687,C535V1783,end_cn535);
C536:CNPU7_7 port map (start_cn,clk,rst,V390C536,V576C536,V714C536,V1095C536,V1208C536,V1688C536,V1784C536,C536V390,C536V576,C536V714,C536V1095,C536V1208,C536V1688,C536V1784,end_cn536);
C537:CNPU7_7 port map (start_cn,clk,rst,V391C537,V481C537,V715C537,V1096C537,V1209C537,V1689C537,V1785C537,C537V391,C537V481,C537V715,C537V1096,C537V1209,C537V1689,C537V1785,end_cn537);
C538:CNPU7_7 port map (start_cn,clk,rst,V392C538,V482C538,V716C538,V1097C538,V1210C538,V1690C538,V1786C538,C538V392,C538V482,C538V716,C538V1097,C538V1210,C538V1690,C538V1786,end_cn538);
C539:CNPU7_7 port map (start_cn,clk,rst,V393C539,V483C539,V717C539,V1098C539,V1211C539,V1691C539,V1787C539,C539V393,C539V483,C539V717,C539V1098,C539V1211,C539V1691,C539V1787,end_cn539);
C540:CNPU7_7 port map (start_cn,clk,rst,V394C540,V484C540,V718C540,V1099C540,V1212C540,V1692C540,V1788C540,C540V394,C540V484,C540V718,C540V1099,C540V1212,C540V1692,C540V1788,end_cn540);
C541:CNPU7_7 port map (start_cn,clk,rst,V395C541,V485C541,V719C541,V1100C541,V1213C541,V1693C541,V1789C541,C541V395,C541V485,C541V719,C541V1100,C541V1213,C541V1693,C541V1789,end_cn541);
C542:CNPU7_7 port map (start_cn,clk,rst,V396C542,V486C542,V720C542,V1101C542,V1214C542,V1694C542,V1790C542,C542V396,C542V486,C542V720,C542V1101,C542V1214,C542V1694,C542V1790,end_cn542);
C543:CNPU7_7 port map (start_cn,clk,rst,V397C543,V487C543,V721C543,V1102C543,V1215C543,V1695C543,V1791C543,C543V397,C543V487,C543V721,C543V1102,C543V1215,C543V1695,C543V1791,end_cn543);
C544:CNPU7_7 port map (start_cn,clk,rst,V398C544,V488C544,V722C544,V1103C544,V1216C544,V1696C544,V1792C544,C544V398,C544V488,C544V722,C544V1103,C544V1216,C544V1696,C544V1792,end_cn544);
C545:CNPU7_7 port map (start_cn,clk,rst,V399C545,V489C545,V723C545,V1104C545,V1217C545,V1697C545,V1793C545,C545V399,C545V489,C545V723,C545V1104,C545V1217,C545V1697,C545V1793,end_cn545);
C546:CNPU7_7 port map (start_cn,clk,rst,V400C546,V490C546,V724C546,V1105C546,V1218C546,V1698C546,V1794C546,C546V400,C546V490,C546V724,C546V1105,C546V1218,C546V1698,C546V1794,end_cn546);
C547:CNPU7_7 port map (start_cn,clk,rst,V401C547,V491C547,V725C547,V1106C547,V1219C547,V1699C547,V1795C547,C547V401,C547V491,C547V725,C547V1106,C547V1219,C547V1699,C547V1795,end_cn547);
C548:CNPU7_7 port map (start_cn,clk,rst,V402C548,V492C548,V726C548,V1107C548,V1220C548,V1700C548,V1796C548,C548V402,C548V492,C548V726,C548V1107,C548V1220,C548V1700,C548V1796,end_cn548);
C549:CNPU7_7 port map (start_cn,clk,rst,V403C549,V493C549,V727C549,V1108C549,V1221C549,V1701C549,V1797C549,C549V403,C549V493,C549V727,C549V1108,C549V1221,C549V1701,C549V1797,end_cn549);
C550:CNPU7_7 port map (start_cn,clk,rst,V404C550,V494C550,V728C550,V1109C550,V1222C550,V1702C550,V1798C550,C550V404,C550V494,C550V728,C550V1109,C550V1222,C550V1702,C550V1798,end_cn550);
C551:CNPU7_7 port map (start_cn,clk,rst,V405C551,V495C551,V729C551,V1110C551,V1223C551,V1703C551,V1799C551,C551V405,C551V495,C551V729,C551V1110,C551V1223,C551V1703,C551V1799,end_cn551);
C552:CNPU7_7 port map (start_cn,clk,rst,V406C552,V496C552,V730C552,V1111C552,V1224C552,V1704C552,V1800C552,C552V406,C552V496,C552V730,C552V1111,C552V1224,C552V1704,C552V1800,end_cn552);
C553:CNPU7_7 port map (start_cn,clk,rst,V407C553,V497C553,V731C553,V1112C553,V1225C553,V1705C553,V1801C553,C553V407,C553V497,C553V731,C553V1112,C553V1225,C553V1705,C553V1801,end_cn553);
C554:CNPU7_7 port map (start_cn,clk,rst,V408C554,V498C554,V732C554,V1113C554,V1226C554,V1706C554,V1802C554,C554V408,C554V498,C554V732,C554V1113,C554V1226,C554V1706,C554V1802,end_cn554);
C555:CNPU7_7 port map (start_cn,clk,rst,V409C555,V499C555,V733C555,V1114C555,V1227C555,V1707C555,V1803C555,C555V409,C555V499,C555V733,C555V1114,C555V1227,C555V1707,C555V1803,end_cn555);
C556:CNPU7_7 port map (start_cn,clk,rst,V410C556,V500C556,V734C556,V1115C556,V1228C556,V1708C556,V1804C556,C556V410,C556V500,C556V734,C556V1115,C556V1228,C556V1708,C556V1804,end_cn556);
C557:CNPU7_7 port map (start_cn,clk,rst,V411C557,V501C557,V735C557,V1116C557,V1229C557,V1709C557,V1805C557,C557V411,C557V501,C557V735,C557V1116,C557V1229,C557V1709,C557V1805,end_cn557);
C558:CNPU7_7 port map (start_cn,clk,rst,V412C558,V502C558,V736C558,V1117C558,V1230C558,V1710C558,V1806C558,C558V412,C558V502,C558V736,C558V1117,C558V1230,C558V1710,C558V1806,end_cn558);
C559:CNPU7_7 port map (start_cn,clk,rst,V413C559,V503C559,V737C559,V1118C559,V1231C559,V1711C559,V1807C559,C559V413,C559V503,C559V737,C559V1118,C559V1231,C559V1711,C559V1807,end_cn559);
C560:CNPU7_7 port map (start_cn,clk,rst,V414C560,V504C560,V738C560,V1119C560,V1232C560,V1712C560,V1808C560,C560V414,C560V504,C560V738,C560V1119,C560V1232,C560V1712,C560V1808,end_cn560);
C561:CNPU7_7 port map (start_cn,clk,rst,V415C561,V505C561,V739C561,V1120C561,V1233C561,V1713C561,V1809C561,C561V415,C561V505,C561V739,C561V1120,C561V1233,C561V1713,C561V1809,end_cn561);
C562:CNPU7_7 port map (start_cn,clk,rst,V416C562,V506C562,V740C562,V1121C562,V1234C562,V1714C562,V1810C562,C562V416,C562V506,C562V740,C562V1121,C562V1234,C562V1714,C562V1810,end_cn562);
C563:CNPU7_7 port map (start_cn,clk,rst,V417C563,V507C563,V741C563,V1122C563,V1235C563,V1715C563,V1811C563,C563V417,C563V507,C563V741,C563V1122,C563V1235,C563V1715,C563V1811,end_cn563);
C564:CNPU7_7 port map (start_cn,clk,rst,V418C564,V508C564,V742C564,V1123C564,V1236C564,V1716C564,V1812C564,C564V418,C564V508,C564V742,C564V1123,C564V1236,C564V1716,C564V1812,end_cn564);
C565:CNPU7_7 port map (start_cn,clk,rst,V419C565,V509C565,V743C565,V1124C565,V1237C565,V1717C565,V1813C565,C565V419,C565V509,C565V743,C565V1124,C565V1237,C565V1717,C565V1813,end_cn565);
C566:CNPU7_7 port map (start_cn,clk,rst,V420C566,V510C566,V744C566,V1125C566,V1238C566,V1718C566,V1814C566,C566V420,C566V510,C566V744,C566V1125,C566V1238,C566V1718,C566V1814,end_cn566);
C567:CNPU7_7 port map (start_cn,clk,rst,V421C567,V511C567,V745C567,V1126C567,V1239C567,V1719C567,V1815C567,C567V421,C567V511,C567V745,C567V1126,C567V1239,C567V1719,C567V1815,end_cn567);
C568:CNPU7_7 port map (start_cn,clk,rst,V422C568,V512C568,V746C568,V1127C568,V1240C568,V1720C568,V1816C568,C568V422,C568V512,C568V746,C568V1127,C568V1240,C568V1720,C568V1816,end_cn568);
C569:CNPU7_7 port map (start_cn,clk,rst,V423C569,V513C569,V747C569,V1128C569,V1241C569,V1721C569,V1817C569,C569V423,C569V513,C569V747,C569V1128,C569V1241,C569V1721,C569V1817,end_cn569);
C570:CNPU7_7 port map (start_cn,clk,rst,V424C570,V514C570,V748C570,V1129C570,V1242C570,V1722C570,V1818C570,C570V424,C570V514,C570V748,C570V1129,C570V1242,C570V1722,C570V1818,end_cn570);
C571:CNPU7_7 port map (start_cn,clk,rst,V425C571,V515C571,V749C571,V1130C571,V1243C571,V1723C571,V1819C571,C571V425,C571V515,C571V749,C571V1130,C571V1243,C571V1723,C571V1819,end_cn571);
C572:CNPU7_7 port map (start_cn,clk,rst,V426C572,V516C572,V750C572,V1131C572,V1244C572,V1724C572,V1820C572,C572V426,C572V516,C572V750,C572V1131,C572V1244,C572V1724,C572V1820,end_cn572);
C573:CNPU7_7 port map (start_cn,clk,rst,V427C573,V517C573,V751C573,V1132C573,V1245C573,V1725C573,V1821C573,C573V427,C573V517,C573V751,C573V1132,C573V1245,C573V1725,C573V1821,end_cn573);
C574:CNPU7_7 port map (start_cn,clk,rst,V428C574,V518C574,V752C574,V1133C574,V1246C574,V1726C574,V1822C574,C574V428,C574V518,C574V752,C574V1133,C574V1246,C574V1726,C574V1822,end_cn574);
C575:CNPU7_7 port map (start_cn,clk,rst,V429C575,V519C575,V753C575,V1134C575,V1247C575,V1727C575,V1823C575,C575V429,C575V519,C575V753,C575V1134,C575V1247,C575V1727,C575V1823,end_cn575);
C576:CNPU7_7 port map (start_cn,clk,rst,V430C576,V520C576,V754C576,V1135C576,V1248C576,V1728C576,V1824C576,C576V430,C576V520,C576V754,C576V1135,C576V1248,C576V1728,C576V1824,end_cn576);
C577:CNPU6_6 port map (start_cn,clk,rst,V288C577,V342C577,V879C577,V979C577,V1729C577,V1825C577,C577V288,C577V342,C577V879,C577V979,C577V1729,C577V1825,end_cn577);
C578:CNPU6_6 port map (start_cn,clk,rst,V193C578,V343C578,V880C578,V980C578,V1730C578,V1826C578,C578V193,C578V343,C578V880,C578V980,C578V1730,C578V1826,end_cn578);
C579:CNPU6_6 port map (start_cn,clk,rst,V194C579,V344C579,V881C579,V981C579,V1731C579,V1827C579,C579V194,C579V344,C579V881,C579V981,C579V1731,C579V1827,end_cn579);
C580:CNPU6_6 port map (start_cn,clk,rst,V195C580,V345C580,V882C580,V982C580,V1732C580,V1828C580,C580V195,C580V345,C580V882,C580V982,C580V1732,C580V1828,end_cn580);
C581:CNPU6_6 port map (start_cn,clk,rst,V196C581,V346C581,V883C581,V983C581,V1733C581,V1829C581,C581V196,C581V346,C581V883,C581V983,C581V1733,C581V1829,end_cn581);
C582:CNPU6_6 port map (start_cn,clk,rst,V197C582,V347C582,V884C582,V984C582,V1734C582,V1830C582,C582V197,C582V347,C582V884,C582V984,C582V1734,C582V1830,end_cn582);
C583:CNPU6_6 port map (start_cn,clk,rst,V198C583,V348C583,V885C583,V985C583,V1735C583,V1831C583,C583V198,C583V348,C583V885,C583V985,C583V1735,C583V1831,end_cn583);
C584:CNPU6_6 port map (start_cn,clk,rst,V199C584,V349C584,V886C584,V986C584,V1736C584,V1832C584,C584V199,C584V349,C584V886,C584V986,C584V1736,C584V1832,end_cn584);
C585:CNPU6_6 port map (start_cn,clk,rst,V200C585,V350C585,V887C585,V987C585,V1737C585,V1833C585,C585V200,C585V350,C585V887,C585V987,C585V1737,C585V1833,end_cn585);
C586:CNPU6_6 port map (start_cn,clk,rst,V201C586,V351C586,V888C586,V988C586,V1738C586,V1834C586,C586V201,C586V351,C586V888,C586V988,C586V1738,C586V1834,end_cn586);
C587:CNPU6_6 port map (start_cn,clk,rst,V202C587,V352C587,V889C587,V989C587,V1739C587,V1835C587,C587V202,C587V352,C587V889,C587V989,C587V1739,C587V1835,end_cn587);
C588:CNPU6_6 port map (start_cn,clk,rst,V203C588,V353C588,V890C588,V990C588,V1740C588,V1836C588,C588V203,C588V353,C588V890,C588V990,C588V1740,C588V1836,end_cn588);
C589:CNPU6_6 port map (start_cn,clk,rst,V204C589,V354C589,V891C589,V991C589,V1741C589,V1837C589,C589V204,C589V354,C589V891,C589V991,C589V1741,C589V1837,end_cn589);
C590:CNPU6_6 port map (start_cn,clk,rst,V205C590,V355C590,V892C590,V992C590,V1742C590,V1838C590,C590V205,C590V355,C590V892,C590V992,C590V1742,C590V1838,end_cn590);
C591:CNPU6_6 port map (start_cn,clk,rst,V206C591,V356C591,V893C591,V993C591,V1743C591,V1839C591,C591V206,C591V356,C591V893,C591V993,C591V1743,C591V1839,end_cn591);
C592:CNPU6_6 port map (start_cn,clk,rst,V207C592,V357C592,V894C592,V994C592,V1744C592,V1840C592,C592V207,C592V357,C592V894,C592V994,C592V1744,C592V1840,end_cn592);
C593:CNPU6_6 port map (start_cn,clk,rst,V208C593,V358C593,V895C593,V995C593,V1745C593,V1841C593,C593V208,C593V358,C593V895,C593V995,C593V1745,C593V1841,end_cn593);
C594:CNPU6_6 port map (start_cn,clk,rst,V209C594,V359C594,V896C594,V996C594,V1746C594,V1842C594,C594V209,C594V359,C594V896,C594V996,C594V1746,C594V1842,end_cn594);
C595:CNPU6_6 port map (start_cn,clk,rst,V210C595,V360C595,V897C595,V997C595,V1747C595,V1843C595,C595V210,C595V360,C595V897,C595V997,C595V1747,C595V1843,end_cn595);
C596:CNPU6_6 port map (start_cn,clk,rst,V211C596,V361C596,V898C596,V998C596,V1748C596,V1844C596,C596V211,C596V361,C596V898,C596V998,C596V1748,C596V1844,end_cn596);
C597:CNPU6_6 port map (start_cn,clk,rst,V212C597,V362C597,V899C597,V999C597,V1749C597,V1845C597,C597V212,C597V362,C597V899,C597V999,C597V1749,C597V1845,end_cn597);
C598:CNPU6_6 port map (start_cn,clk,rst,V213C598,V363C598,V900C598,V1000C598,V1750C598,V1846C598,C598V213,C598V363,C598V900,C598V1000,C598V1750,C598V1846,end_cn598);
C599:CNPU6_6 port map (start_cn,clk,rst,V214C599,V364C599,V901C599,V1001C599,V1751C599,V1847C599,C599V214,C599V364,C599V901,C599V1001,C599V1751,C599V1847,end_cn599);
C600:CNPU6_6 port map (start_cn,clk,rst,V215C600,V365C600,V902C600,V1002C600,V1752C600,V1848C600,C600V215,C600V365,C600V902,C600V1002,C600V1752,C600V1848,end_cn600);
C601:CNPU6_6 port map (start_cn,clk,rst,V216C601,V366C601,V903C601,V1003C601,V1753C601,V1849C601,C601V216,C601V366,C601V903,C601V1003,C601V1753,C601V1849,end_cn601);
C602:CNPU6_6 port map (start_cn,clk,rst,V217C602,V367C602,V904C602,V1004C602,V1754C602,V1850C602,C602V217,C602V367,C602V904,C602V1004,C602V1754,C602V1850,end_cn602);
C603:CNPU6_6 port map (start_cn,clk,rst,V218C603,V368C603,V905C603,V1005C603,V1755C603,V1851C603,C603V218,C603V368,C603V905,C603V1005,C603V1755,C603V1851,end_cn603);
C604:CNPU6_6 port map (start_cn,clk,rst,V219C604,V369C604,V906C604,V1006C604,V1756C604,V1852C604,C604V219,C604V369,C604V906,C604V1006,C604V1756,C604V1852,end_cn604);
C605:CNPU6_6 port map (start_cn,clk,rst,V220C605,V370C605,V907C605,V1007C605,V1757C605,V1853C605,C605V220,C605V370,C605V907,C605V1007,C605V1757,C605V1853,end_cn605);
C606:CNPU6_6 port map (start_cn,clk,rst,V221C606,V371C606,V908C606,V1008C606,V1758C606,V1854C606,C606V221,C606V371,C606V908,C606V1008,C606V1758,C606V1854,end_cn606);
C607:CNPU6_6 port map (start_cn,clk,rst,V222C607,V372C607,V909C607,V1009C607,V1759C607,V1855C607,C607V222,C607V372,C607V909,C607V1009,C607V1759,C607V1855,end_cn607);
C608:CNPU6_6 port map (start_cn,clk,rst,V223C608,V373C608,V910C608,V1010C608,V1760C608,V1856C608,C608V223,C608V373,C608V910,C608V1010,C608V1760,C608V1856,end_cn608);
C609:CNPU6_6 port map (start_cn,clk,rst,V224C609,V374C609,V911C609,V1011C609,V1761C609,V1857C609,C609V224,C609V374,C609V911,C609V1011,C609V1761,C609V1857,end_cn609);
C610:CNPU6_6 port map (start_cn,clk,rst,V225C610,V375C610,V912C610,V1012C610,V1762C610,V1858C610,C610V225,C610V375,C610V912,C610V1012,C610V1762,C610V1858,end_cn610);
C611:CNPU6_6 port map (start_cn,clk,rst,V226C611,V376C611,V913C611,V1013C611,V1763C611,V1859C611,C611V226,C611V376,C611V913,C611V1013,C611V1763,C611V1859,end_cn611);
C612:CNPU6_6 port map (start_cn,clk,rst,V227C612,V377C612,V914C612,V1014C612,V1764C612,V1860C612,C612V227,C612V377,C612V914,C612V1014,C612V1764,C612V1860,end_cn612);
C613:CNPU6_6 port map (start_cn,clk,rst,V228C613,V378C613,V915C613,V1015C613,V1765C613,V1861C613,C613V228,C613V378,C613V915,C613V1015,C613V1765,C613V1861,end_cn613);
C614:CNPU6_6 port map (start_cn,clk,rst,V229C614,V379C614,V916C614,V1016C614,V1766C614,V1862C614,C614V229,C614V379,C614V916,C614V1016,C614V1766,C614V1862,end_cn614);
C615:CNPU6_6 port map (start_cn,clk,rst,V230C615,V380C615,V917C615,V1017C615,V1767C615,V1863C615,C615V230,C615V380,C615V917,C615V1017,C615V1767,C615V1863,end_cn615);
C616:CNPU6_6 port map (start_cn,clk,rst,V231C616,V381C616,V918C616,V1018C616,V1768C616,V1864C616,C616V231,C616V381,C616V918,C616V1018,C616V1768,C616V1864,end_cn616);
C617:CNPU6_6 port map (start_cn,clk,rst,V232C617,V382C617,V919C617,V1019C617,V1769C617,V1865C617,C617V232,C617V382,C617V919,C617V1019,C617V1769,C617V1865,end_cn617);
C618:CNPU6_6 port map (start_cn,clk,rst,V233C618,V383C618,V920C618,V1020C618,V1770C618,V1866C618,C618V233,C618V383,C618V920,C618V1020,C618V1770,C618V1866,end_cn618);
C619:CNPU6_6 port map (start_cn,clk,rst,V234C619,V384C619,V921C619,V1021C619,V1771C619,V1867C619,C619V234,C619V384,C619V921,C619V1021,C619V1771,C619V1867,end_cn619);
C620:CNPU6_6 port map (start_cn,clk,rst,V235C620,V289C620,V922C620,V1022C620,V1772C620,V1868C620,C620V235,C620V289,C620V922,C620V1022,C620V1772,C620V1868,end_cn620);
C621:CNPU6_6 port map (start_cn,clk,rst,V236C621,V290C621,V923C621,V1023C621,V1773C621,V1869C621,C621V236,C621V290,C621V923,C621V1023,C621V1773,C621V1869,end_cn621);
C622:CNPU6_6 port map (start_cn,clk,rst,V237C622,V291C622,V924C622,V1024C622,V1774C622,V1870C622,C622V237,C622V291,C622V924,C622V1024,C622V1774,C622V1870,end_cn622);
C623:CNPU6_6 port map (start_cn,clk,rst,V238C623,V292C623,V925C623,V1025C623,V1775C623,V1871C623,C623V238,C623V292,C623V925,C623V1025,C623V1775,C623V1871,end_cn623);
C624:CNPU6_6 port map (start_cn,clk,rst,V239C624,V293C624,V926C624,V1026C624,V1776C624,V1872C624,C624V239,C624V293,C624V926,C624V1026,C624V1776,C624V1872,end_cn624);
C625:CNPU6_6 port map (start_cn,clk,rst,V240C625,V294C625,V927C625,V1027C625,V1777C625,V1873C625,C625V240,C625V294,C625V927,C625V1027,C625V1777,C625V1873,end_cn625);
C626:CNPU6_6 port map (start_cn,clk,rst,V241C626,V295C626,V928C626,V1028C626,V1778C626,V1874C626,C626V241,C626V295,C626V928,C626V1028,C626V1778,C626V1874,end_cn626);
C627:CNPU6_6 port map (start_cn,clk,rst,V242C627,V296C627,V929C627,V1029C627,V1779C627,V1875C627,C627V242,C627V296,C627V929,C627V1029,C627V1779,C627V1875,end_cn627);
C628:CNPU6_6 port map (start_cn,clk,rst,V243C628,V297C628,V930C628,V1030C628,V1780C628,V1876C628,C628V243,C628V297,C628V930,C628V1030,C628V1780,C628V1876,end_cn628);
C629:CNPU6_6 port map (start_cn,clk,rst,V244C629,V298C629,V931C629,V1031C629,V1781C629,V1877C629,C629V244,C629V298,C629V931,C629V1031,C629V1781,C629V1877,end_cn629);
C630:CNPU6_6 port map (start_cn,clk,rst,V245C630,V299C630,V932C630,V1032C630,V1782C630,V1878C630,C630V245,C630V299,C630V932,C630V1032,C630V1782,C630V1878,end_cn630);
C631:CNPU6_6 port map (start_cn,clk,rst,V246C631,V300C631,V933C631,V1033C631,V1783C631,V1879C631,C631V246,C631V300,C631V933,C631V1033,C631V1783,C631V1879,end_cn631);
C632:CNPU6_6 port map (start_cn,clk,rst,V247C632,V301C632,V934C632,V1034C632,V1784C632,V1880C632,C632V247,C632V301,C632V934,C632V1034,C632V1784,C632V1880,end_cn632);
C633:CNPU6_6 port map (start_cn,clk,rst,V248C633,V302C633,V935C633,V1035C633,V1785C633,V1881C633,C633V248,C633V302,C633V935,C633V1035,C633V1785,C633V1881,end_cn633);
C634:CNPU6_6 port map (start_cn,clk,rst,V249C634,V303C634,V936C634,V1036C634,V1786C634,V1882C634,C634V249,C634V303,C634V936,C634V1036,C634V1786,C634V1882,end_cn634);
C635:CNPU6_6 port map (start_cn,clk,rst,V250C635,V304C635,V937C635,V1037C635,V1787C635,V1883C635,C635V250,C635V304,C635V937,C635V1037,C635V1787,C635V1883,end_cn635);
C636:CNPU6_6 port map (start_cn,clk,rst,V251C636,V305C636,V938C636,V1038C636,V1788C636,V1884C636,C636V251,C636V305,C636V938,C636V1038,C636V1788,C636V1884,end_cn636);
C637:CNPU6_6 port map (start_cn,clk,rst,V252C637,V306C637,V939C637,V1039C637,V1789C637,V1885C637,C637V252,C637V306,C637V939,C637V1039,C637V1789,C637V1885,end_cn637);
C638:CNPU6_6 port map (start_cn,clk,rst,V253C638,V307C638,V940C638,V1040C638,V1790C638,V1886C638,C638V253,C638V307,C638V940,C638V1040,C638V1790,C638V1886,end_cn638);
C639:CNPU6_6 port map (start_cn,clk,rst,V254C639,V308C639,V941C639,V1041C639,V1791C639,V1887C639,C639V254,C639V308,C639V941,C639V1041,C639V1791,C639V1887,end_cn639);
C640:CNPU6_6 port map (start_cn,clk,rst,V255C640,V309C640,V942C640,V1042C640,V1792C640,V1888C640,C640V255,C640V309,C640V942,C640V1042,C640V1792,C640V1888,end_cn640);
C641:CNPU6_6 port map (start_cn,clk,rst,V256C641,V310C641,V943C641,V1043C641,V1793C641,V1889C641,C641V256,C641V310,C641V943,C641V1043,C641V1793,C641V1889,end_cn641);
C642:CNPU6_6 port map (start_cn,clk,rst,V257C642,V311C642,V944C642,V1044C642,V1794C642,V1890C642,C642V257,C642V311,C642V944,C642V1044,C642V1794,C642V1890,end_cn642);
C643:CNPU6_6 port map (start_cn,clk,rst,V258C643,V312C643,V945C643,V1045C643,V1795C643,V1891C643,C643V258,C643V312,C643V945,C643V1045,C643V1795,C643V1891,end_cn643);
C644:CNPU6_6 port map (start_cn,clk,rst,V259C644,V313C644,V946C644,V1046C644,V1796C644,V1892C644,C644V259,C644V313,C644V946,C644V1046,C644V1796,C644V1892,end_cn644);
C645:CNPU6_6 port map (start_cn,clk,rst,V260C645,V314C645,V947C645,V1047C645,V1797C645,V1893C645,C645V260,C645V314,C645V947,C645V1047,C645V1797,C645V1893,end_cn645);
C646:CNPU6_6 port map (start_cn,clk,rst,V261C646,V315C646,V948C646,V1048C646,V1798C646,V1894C646,C646V261,C646V315,C646V948,C646V1048,C646V1798,C646V1894,end_cn646);
C647:CNPU6_6 port map (start_cn,clk,rst,V262C647,V316C647,V949C647,V1049C647,V1799C647,V1895C647,C647V262,C647V316,C647V949,C647V1049,C647V1799,C647V1895,end_cn647);
C648:CNPU6_6 port map (start_cn,clk,rst,V263C648,V317C648,V950C648,V1050C648,V1800C648,V1896C648,C648V263,C648V317,C648V950,C648V1050,C648V1800,C648V1896,end_cn648);
C649:CNPU6_6 port map (start_cn,clk,rst,V264C649,V318C649,V951C649,V1051C649,V1801C649,V1897C649,C649V264,C649V318,C649V951,C649V1051,C649V1801,C649V1897,end_cn649);
C650:CNPU6_6 port map (start_cn,clk,rst,V265C650,V319C650,V952C650,V1052C650,V1802C650,V1898C650,C650V265,C650V319,C650V952,C650V1052,C650V1802,C650V1898,end_cn650);
C651:CNPU6_6 port map (start_cn,clk,rst,V266C651,V320C651,V953C651,V1053C651,V1803C651,V1899C651,C651V266,C651V320,C651V953,C651V1053,C651V1803,C651V1899,end_cn651);
C652:CNPU6_6 port map (start_cn,clk,rst,V267C652,V321C652,V954C652,V1054C652,V1804C652,V1900C652,C652V267,C652V321,C652V954,C652V1054,C652V1804,C652V1900,end_cn652);
C653:CNPU6_6 port map (start_cn,clk,rst,V268C653,V322C653,V955C653,V1055C653,V1805C653,V1901C653,C653V268,C653V322,C653V955,C653V1055,C653V1805,C653V1901,end_cn653);
C654:CNPU6_6 port map (start_cn,clk,rst,V269C654,V323C654,V956C654,V1056C654,V1806C654,V1902C654,C654V269,C654V323,C654V956,C654V1056,C654V1806,C654V1902,end_cn654);
C655:CNPU6_6 port map (start_cn,clk,rst,V270C655,V324C655,V957C655,V961C655,V1807C655,V1903C655,C655V270,C655V324,C655V957,C655V961,C655V1807,C655V1903,end_cn655);
C656:CNPU6_6 port map (start_cn,clk,rst,V271C656,V325C656,V958C656,V962C656,V1808C656,V1904C656,C656V271,C656V325,C656V958,C656V962,C656V1808,C656V1904,end_cn656);
C657:CNPU6_6 port map (start_cn,clk,rst,V272C657,V326C657,V959C657,V963C657,V1809C657,V1905C657,C657V272,C657V326,C657V959,C657V963,C657V1809,C657V1905,end_cn657);
C658:CNPU6_6 port map (start_cn,clk,rst,V273C658,V327C658,V960C658,V964C658,V1810C658,V1906C658,C658V273,C658V327,C658V960,C658V964,C658V1810,C658V1906,end_cn658);
C659:CNPU6_6 port map (start_cn,clk,rst,V274C659,V328C659,V865C659,V965C659,V1811C659,V1907C659,C659V274,C659V328,C659V865,C659V965,C659V1811,C659V1907,end_cn659);
C660:CNPU6_6 port map (start_cn,clk,rst,V275C660,V329C660,V866C660,V966C660,V1812C660,V1908C660,C660V275,C660V329,C660V866,C660V966,C660V1812,C660V1908,end_cn660);
C661:CNPU6_6 port map (start_cn,clk,rst,V276C661,V330C661,V867C661,V967C661,V1813C661,V1909C661,C661V276,C661V330,C661V867,C661V967,C661V1813,C661V1909,end_cn661);
C662:CNPU6_6 port map (start_cn,clk,rst,V277C662,V331C662,V868C662,V968C662,V1814C662,V1910C662,C662V277,C662V331,C662V868,C662V968,C662V1814,C662V1910,end_cn662);
C663:CNPU6_6 port map (start_cn,clk,rst,V278C663,V332C663,V869C663,V969C663,V1815C663,V1911C663,C663V278,C663V332,C663V869,C663V969,C663V1815,C663V1911,end_cn663);
C664:CNPU6_6 port map (start_cn,clk,rst,V279C664,V333C664,V870C664,V970C664,V1816C664,V1912C664,C664V279,C664V333,C664V870,C664V970,C664V1816,C664V1912,end_cn664);
C665:CNPU6_6 port map (start_cn,clk,rst,V280C665,V334C665,V871C665,V971C665,V1817C665,V1913C665,C665V280,C665V334,C665V871,C665V971,C665V1817,C665V1913,end_cn665);
C666:CNPU6_6 port map (start_cn,clk,rst,V281C666,V335C666,V872C666,V972C666,V1818C666,V1914C666,C666V281,C666V335,C666V872,C666V972,C666V1818,C666V1914,end_cn666);
C667:CNPU6_6 port map (start_cn,clk,rst,V282C667,V336C667,V873C667,V973C667,V1819C667,V1915C667,C667V282,C667V336,C667V873,C667V973,C667V1819,C667V1915,end_cn667);
C668:CNPU6_6 port map (start_cn,clk,rst,V283C668,V337C668,V874C668,V974C668,V1820C668,V1916C668,C668V283,C668V337,C668V874,C668V974,C668V1820,C668V1916,end_cn668);
C669:CNPU6_6 port map (start_cn,clk,rst,V284C669,V338C669,V875C669,V975C669,V1821C669,V1917C669,C669V284,C669V338,C669V875,C669V975,C669V1821,C669V1917,end_cn669);
C670:CNPU6_6 port map (start_cn,clk,rst,V285C670,V339C670,V876C670,V976C670,V1822C670,V1918C670,C670V285,C670V339,C670V876,C670V976,C670V1822,C670V1918,end_cn670);
C671:CNPU6_6 port map (start_cn,clk,rst,V286C671,V340C671,V877C671,V977C671,V1823C671,V1919C671,C671V286,C671V340,C671V877,C671V977,C671V1823,C671V1919,end_cn671);
C672:CNPU6_6 port map (start_cn,clk,rst,V287C672,V341C672,V878C672,V978C672,V1824C672,V1920C672,C672V287,C672V341,C672V878,C672V978,C672V1824,C672V1920,end_cn672);
C673:CNPU6_6 port map (start_cn,clk,rst,V108C673,V266C673,V579C673,V912C673,V1825C673,V1921C673,C673V108,C673V266,C673V579,C673V912,C673V1825,C673V1921,end_cn673);
C674:CNPU6_6 port map (start_cn,clk,rst,V109C674,V267C674,V580C674,V913C674,V1826C674,V1922C674,C674V109,C674V267,C674V580,C674V913,C674V1826,C674V1922,end_cn674);
C675:CNPU6_6 port map (start_cn,clk,rst,V110C675,V268C675,V581C675,V914C675,V1827C675,V1923C675,C675V110,C675V268,C675V581,C675V914,C675V1827,C675V1923,end_cn675);
C676:CNPU6_6 port map (start_cn,clk,rst,V111C676,V269C676,V582C676,V915C676,V1828C676,V1924C676,C676V111,C676V269,C676V582,C676V915,C676V1828,C676V1924,end_cn676);
C677:CNPU6_6 port map (start_cn,clk,rst,V112C677,V270C677,V583C677,V916C677,V1829C677,V1925C677,C677V112,C677V270,C677V583,C677V916,C677V1829,C677V1925,end_cn677);
C678:CNPU6_6 port map (start_cn,clk,rst,V113C678,V271C678,V584C678,V917C678,V1830C678,V1926C678,C678V113,C678V271,C678V584,C678V917,C678V1830,C678V1926,end_cn678);
C679:CNPU6_6 port map (start_cn,clk,rst,V114C679,V272C679,V585C679,V918C679,V1831C679,V1927C679,C679V114,C679V272,C679V585,C679V918,C679V1831,C679V1927,end_cn679);
C680:CNPU6_6 port map (start_cn,clk,rst,V115C680,V273C680,V586C680,V919C680,V1832C680,V1928C680,C680V115,C680V273,C680V586,C680V919,C680V1832,C680V1928,end_cn680);
C681:CNPU6_6 port map (start_cn,clk,rst,V116C681,V274C681,V587C681,V920C681,V1833C681,V1929C681,C681V116,C681V274,C681V587,C681V920,C681V1833,C681V1929,end_cn681);
C682:CNPU6_6 port map (start_cn,clk,rst,V117C682,V275C682,V588C682,V921C682,V1834C682,V1930C682,C682V117,C682V275,C682V588,C682V921,C682V1834,C682V1930,end_cn682);
C683:CNPU6_6 port map (start_cn,clk,rst,V118C683,V276C683,V589C683,V922C683,V1835C683,V1931C683,C683V118,C683V276,C683V589,C683V922,C683V1835,C683V1931,end_cn683);
C684:CNPU6_6 port map (start_cn,clk,rst,V119C684,V277C684,V590C684,V923C684,V1836C684,V1932C684,C684V119,C684V277,C684V590,C684V923,C684V1836,C684V1932,end_cn684);
C685:CNPU6_6 port map (start_cn,clk,rst,V120C685,V278C685,V591C685,V924C685,V1837C685,V1933C685,C685V120,C685V278,C685V591,C685V924,C685V1837,C685V1933,end_cn685);
C686:CNPU6_6 port map (start_cn,clk,rst,V121C686,V279C686,V592C686,V925C686,V1838C686,V1934C686,C686V121,C686V279,C686V592,C686V925,C686V1838,C686V1934,end_cn686);
C687:CNPU6_6 port map (start_cn,clk,rst,V122C687,V280C687,V593C687,V926C687,V1839C687,V1935C687,C687V122,C687V280,C687V593,C687V926,C687V1839,C687V1935,end_cn687);
C688:CNPU6_6 port map (start_cn,clk,rst,V123C688,V281C688,V594C688,V927C688,V1840C688,V1936C688,C688V123,C688V281,C688V594,C688V927,C688V1840,C688V1936,end_cn688);
C689:CNPU6_6 port map (start_cn,clk,rst,V124C689,V282C689,V595C689,V928C689,V1841C689,V1937C689,C689V124,C689V282,C689V595,C689V928,C689V1841,C689V1937,end_cn689);
C690:CNPU6_6 port map (start_cn,clk,rst,V125C690,V283C690,V596C690,V929C690,V1842C690,V1938C690,C690V125,C690V283,C690V596,C690V929,C690V1842,C690V1938,end_cn690);
C691:CNPU6_6 port map (start_cn,clk,rst,V126C691,V284C691,V597C691,V930C691,V1843C691,V1939C691,C691V126,C691V284,C691V597,C691V930,C691V1843,C691V1939,end_cn691);
C692:CNPU6_6 port map (start_cn,clk,rst,V127C692,V285C692,V598C692,V931C692,V1844C692,V1940C692,C692V127,C692V285,C692V598,C692V931,C692V1844,C692V1940,end_cn692);
C693:CNPU6_6 port map (start_cn,clk,rst,V128C693,V286C693,V599C693,V932C693,V1845C693,V1941C693,C693V128,C693V286,C693V599,C693V932,C693V1845,C693V1941,end_cn693);
C694:CNPU6_6 port map (start_cn,clk,rst,V129C694,V287C694,V600C694,V933C694,V1846C694,V1942C694,C694V129,C694V287,C694V600,C694V933,C694V1846,C694V1942,end_cn694);
C695:CNPU6_6 port map (start_cn,clk,rst,V130C695,V288C695,V601C695,V934C695,V1847C695,V1943C695,C695V130,C695V288,C695V601,C695V934,C695V1847,C695V1943,end_cn695);
C696:CNPU6_6 port map (start_cn,clk,rst,V131C696,V193C696,V602C696,V935C696,V1848C696,V1944C696,C696V131,C696V193,C696V602,C696V935,C696V1848,C696V1944,end_cn696);
C697:CNPU6_6 port map (start_cn,clk,rst,V132C697,V194C697,V603C697,V936C697,V1849C697,V1945C697,C697V132,C697V194,C697V603,C697V936,C697V1849,C697V1945,end_cn697);
C698:CNPU6_6 port map (start_cn,clk,rst,V133C698,V195C698,V604C698,V937C698,V1850C698,V1946C698,C698V133,C698V195,C698V604,C698V937,C698V1850,C698V1946,end_cn698);
C699:CNPU6_6 port map (start_cn,clk,rst,V134C699,V196C699,V605C699,V938C699,V1851C699,V1947C699,C699V134,C699V196,C699V605,C699V938,C699V1851,C699V1947,end_cn699);
C700:CNPU6_6 port map (start_cn,clk,rst,V135C700,V197C700,V606C700,V939C700,V1852C700,V1948C700,C700V135,C700V197,C700V606,C700V939,C700V1852,C700V1948,end_cn700);
C701:CNPU6_6 port map (start_cn,clk,rst,V136C701,V198C701,V607C701,V940C701,V1853C701,V1949C701,C701V136,C701V198,C701V607,C701V940,C701V1853,C701V1949,end_cn701);
C702:CNPU6_6 port map (start_cn,clk,rst,V137C702,V199C702,V608C702,V941C702,V1854C702,V1950C702,C702V137,C702V199,C702V608,C702V941,C702V1854,C702V1950,end_cn702);
C703:CNPU6_6 port map (start_cn,clk,rst,V138C703,V200C703,V609C703,V942C703,V1855C703,V1951C703,C703V138,C703V200,C703V609,C703V942,C703V1855,C703V1951,end_cn703);
C704:CNPU6_6 port map (start_cn,clk,rst,V139C704,V201C704,V610C704,V943C704,V1856C704,V1952C704,C704V139,C704V201,C704V610,C704V943,C704V1856,C704V1952,end_cn704);
C705:CNPU6_6 port map (start_cn,clk,rst,V140C705,V202C705,V611C705,V944C705,V1857C705,V1953C705,C705V140,C705V202,C705V611,C705V944,C705V1857,C705V1953,end_cn705);
C706:CNPU6_6 port map (start_cn,clk,rst,V141C706,V203C706,V612C706,V945C706,V1858C706,V1954C706,C706V141,C706V203,C706V612,C706V945,C706V1858,C706V1954,end_cn706);
C707:CNPU6_6 port map (start_cn,clk,rst,V142C707,V204C707,V613C707,V946C707,V1859C707,V1955C707,C707V142,C707V204,C707V613,C707V946,C707V1859,C707V1955,end_cn707);
C708:CNPU6_6 port map (start_cn,clk,rst,V143C708,V205C708,V614C708,V947C708,V1860C708,V1956C708,C708V143,C708V205,C708V614,C708V947,C708V1860,C708V1956,end_cn708);
C709:CNPU6_6 port map (start_cn,clk,rst,V144C709,V206C709,V615C709,V948C709,V1861C709,V1957C709,C709V144,C709V206,C709V615,C709V948,C709V1861,C709V1957,end_cn709);
C710:CNPU6_6 port map (start_cn,clk,rst,V145C710,V207C710,V616C710,V949C710,V1862C710,V1958C710,C710V145,C710V207,C710V616,C710V949,C710V1862,C710V1958,end_cn710);
C711:CNPU6_6 port map (start_cn,clk,rst,V146C711,V208C711,V617C711,V950C711,V1863C711,V1959C711,C711V146,C711V208,C711V617,C711V950,C711V1863,C711V1959,end_cn711);
C712:CNPU6_6 port map (start_cn,clk,rst,V147C712,V209C712,V618C712,V951C712,V1864C712,V1960C712,C712V147,C712V209,C712V618,C712V951,C712V1864,C712V1960,end_cn712);
C713:CNPU6_6 port map (start_cn,clk,rst,V148C713,V210C713,V619C713,V952C713,V1865C713,V1961C713,C713V148,C713V210,C713V619,C713V952,C713V1865,C713V1961,end_cn713);
C714:CNPU6_6 port map (start_cn,clk,rst,V149C714,V211C714,V620C714,V953C714,V1866C714,V1962C714,C714V149,C714V211,C714V620,C714V953,C714V1866,C714V1962,end_cn714);
C715:CNPU6_6 port map (start_cn,clk,rst,V150C715,V212C715,V621C715,V954C715,V1867C715,V1963C715,C715V150,C715V212,C715V621,C715V954,C715V1867,C715V1963,end_cn715);
C716:CNPU6_6 port map (start_cn,clk,rst,V151C716,V213C716,V622C716,V955C716,V1868C716,V1964C716,C716V151,C716V213,C716V622,C716V955,C716V1868,C716V1964,end_cn716);
C717:CNPU6_6 port map (start_cn,clk,rst,V152C717,V214C717,V623C717,V956C717,V1869C717,V1965C717,C717V152,C717V214,C717V623,C717V956,C717V1869,C717V1965,end_cn717);
C718:CNPU6_6 port map (start_cn,clk,rst,V153C718,V215C718,V624C718,V957C718,V1870C718,V1966C718,C718V153,C718V215,C718V624,C718V957,C718V1870,C718V1966,end_cn718);
C719:CNPU6_6 port map (start_cn,clk,rst,V154C719,V216C719,V625C719,V958C719,V1871C719,V1967C719,C719V154,C719V216,C719V625,C719V958,C719V1871,C719V1967,end_cn719);
C720:CNPU6_6 port map (start_cn,clk,rst,V155C720,V217C720,V626C720,V959C720,V1872C720,V1968C720,C720V155,C720V217,C720V626,C720V959,C720V1872,C720V1968,end_cn720);
C721:CNPU6_6 port map (start_cn,clk,rst,V156C721,V218C721,V627C721,V960C721,V1873C721,V1969C721,C721V156,C721V218,C721V627,C721V960,C721V1873,C721V1969,end_cn721);
C722:CNPU6_6 port map (start_cn,clk,rst,V157C722,V219C722,V628C722,V865C722,V1874C722,V1970C722,C722V157,C722V219,C722V628,C722V865,C722V1874,C722V1970,end_cn722);
C723:CNPU6_6 port map (start_cn,clk,rst,V158C723,V220C723,V629C723,V866C723,V1875C723,V1971C723,C723V158,C723V220,C723V629,C723V866,C723V1875,C723V1971,end_cn723);
C724:CNPU6_6 port map (start_cn,clk,rst,V159C724,V221C724,V630C724,V867C724,V1876C724,V1972C724,C724V159,C724V221,C724V630,C724V867,C724V1876,C724V1972,end_cn724);
C725:CNPU6_6 port map (start_cn,clk,rst,V160C725,V222C725,V631C725,V868C725,V1877C725,V1973C725,C725V160,C725V222,C725V631,C725V868,C725V1877,C725V1973,end_cn725);
C726:CNPU6_6 port map (start_cn,clk,rst,V161C726,V223C726,V632C726,V869C726,V1878C726,V1974C726,C726V161,C726V223,C726V632,C726V869,C726V1878,C726V1974,end_cn726);
C727:CNPU6_6 port map (start_cn,clk,rst,V162C727,V224C727,V633C727,V870C727,V1879C727,V1975C727,C727V162,C727V224,C727V633,C727V870,C727V1879,C727V1975,end_cn727);
C728:CNPU6_6 port map (start_cn,clk,rst,V163C728,V225C728,V634C728,V871C728,V1880C728,V1976C728,C728V163,C728V225,C728V634,C728V871,C728V1880,C728V1976,end_cn728);
C729:CNPU6_6 port map (start_cn,clk,rst,V164C729,V226C729,V635C729,V872C729,V1881C729,V1977C729,C729V164,C729V226,C729V635,C729V872,C729V1881,C729V1977,end_cn729);
C730:CNPU6_6 port map (start_cn,clk,rst,V165C730,V227C730,V636C730,V873C730,V1882C730,V1978C730,C730V165,C730V227,C730V636,C730V873,C730V1882,C730V1978,end_cn730);
C731:CNPU6_6 port map (start_cn,clk,rst,V166C731,V228C731,V637C731,V874C731,V1883C731,V1979C731,C731V166,C731V228,C731V637,C731V874,C731V1883,C731V1979,end_cn731);
C732:CNPU6_6 port map (start_cn,clk,rst,V167C732,V229C732,V638C732,V875C732,V1884C732,V1980C732,C732V167,C732V229,C732V638,C732V875,C732V1884,C732V1980,end_cn732);
C733:CNPU6_6 port map (start_cn,clk,rst,V168C733,V230C733,V639C733,V876C733,V1885C733,V1981C733,C733V168,C733V230,C733V639,C733V876,C733V1885,C733V1981,end_cn733);
C734:CNPU6_6 port map (start_cn,clk,rst,V169C734,V231C734,V640C734,V877C734,V1886C734,V1982C734,C734V169,C734V231,C734V640,C734V877,C734V1886,C734V1982,end_cn734);
C735:CNPU6_6 port map (start_cn,clk,rst,V170C735,V232C735,V641C735,V878C735,V1887C735,V1983C735,C735V170,C735V232,C735V641,C735V878,C735V1887,C735V1983,end_cn735);
C736:CNPU6_6 port map (start_cn,clk,rst,V171C736,V233C736,V642C736,V879C736,V1888C736,V1984C736,C736V171,C736V233,C736V642,C736V879,C736V1888,C736V1984,end_cn736);
C737:CNPU6_6 port map (start_cn,clk,rst,V172C737,V234C737,V643C737,V880C737,V1889C737,V1985C737,C737V172,C737V234,C737V643,C737V880,C737V1889,C737V1985,end_cn737);
C738:CNPU6_6 port map (start_cn,clk,rst,V173C738,V235C738,V644C738,V881C738,V1890C738,V1986C738,C738V173,C738V235,C738V644,C738V881,C738V1890,C738V1986,end_cn738);
C739:CNPU6_6 port map (start_cn,clk,rst,V174C739,V236C739,V645C739,V882C739,V1891C739,V1987C739,C739V174,C739V236,C739V645,C739V882,C739V1891,C739V1987,end_cn739);
C740:CNPU6_6 port map (start_cn,clk,rst,V175C740,V237C740,V646C740,V883C740,V1892C740,V1988C740,C740V175,C740V237,C740V646,C740V883,C740V1892,C740V1988,end_cn740);
C741:CNPU6_6 port map (start_cn,clk,rst,V176C741,V238C741,V647C741,V884C741,V1893C741,V1989C741,C741V176,C741V238,C741V647,C741V884,C741V1893,C741V1989,end_cn741);
C742:CNPU6_6 port map (start_cn,clk,rst,V177C742,V239C742,V648C742,V885C742,V1894C742,V1990C742,C742V177,C742V239,C742V648,C742V885,C742V1894,C742V1990,end_cn742);
C743:CNPU6_6 port map (start_cn,clk,rst,V178C743,V240C743,V649C743,V886C743,V1895C743,V1991C743,C743V178,C743V240,C743V649,C743V886,C743V1895,C743V1991,end_cn743);
C744:CNPU6_6 port map (start_cn,clk,rst,V179C744,V241C744,V650C744,V887C744,V1896C744,V1992C744,C744V179,C744V241,C744V650,C744V887,C744V1896,C744V1992,end_cn744);
C745:CNPU6_6 port map (start_cn,clk,rst,V180C745,V242C745,V651C745,V888C745,V1897C745,V1993C745,C745V180,C745V242,C745V651,C745V888,C745V1897,C745V1993,end_cn745);
C746:CNPU6_6 port map (start_cn,clk,rst,V181C746,V243C746,V652C746,V889C746,V1898C746,V1994C746,C746V181,C746V243,C746V652,C746V889,C746V1898,C746V1994,end_cn746);
C747:CNPU6_6 port map (start_cn,clk,rst,V182C747,V244C747,V653C747,V890C747,V1899C747,V1995C747,C747V182,C747V244,C747V653,C747V890,C747V1899,C747V1995,end_cn747);
C748:CNPU6_6 port map (start_cn,clk,rst,V183C748,V245C748,V654C748,V891C748,V1900C748,V1996C748,C748V183,C748V245,C748V654,C748V891,C748V1900,C748V1996,end_cn748);
C749:CNPU6_6 port map (start_cn,clk,rst,V184C749,V246C749,V655C749,V892C749,V1901C749,V1997C749,C749V184,C749V246,C749V655,C749V892,C749V1901,C749V1997,end_cn749);
C750:CNPU6_6 port map (start_cn,clk,rst,V185C750,V247C750,V656C750,V893C750,V1902C750,V1998C750,C750V185,C750V247,C750V656,C750V893,C750V1902,C750V1998,end_cn750);
C751:CNPU6_6 port map (start_cn,clk,rst,V186C751,V248C751,V657C751,V894C751,V1903C751,V1999C751,C751V186,C751V248,C751V657,C751V894,C751V1903,C751V1999,end_cn751);
C752:CNPU6_6 port map (start_cn,clk,rst,V187C752,V249C752,V658C752,V895C752,V1904C752,V2000C752,C752V187,C752V249,C752V658,C752V895,C752V1904,C752V2000,end_cn752);
C753:CNPU6_6 port map (start_cn,clk,rst,V188C753,V250C753,V659C753,V896C753,V1905C753,V2001C753,C753V188,C753V250,C753V659,C753V896,C753V1905,C753V2001,end_cn753);
C754:CNPU6_6 port map (start_cn,clk,rst,V189C754,V251C754,V660C754,V897C754,V1906C754,V2002C754,C754V189,C754V251,C754V660,C754V897,C754V1906,C754V2002,end_cn754);
C755:CNPU6_6 port map (start_cn,clk,rst,V190C755,V252C755,V661C755,V898C755,V1907C755,V2003C755,C755V190,C755V252,C755V661,C755V898,C755V1907,C755V2003,end_cn755);
C756:CNPU6_6 port map (start_cn,clk,rst,V191C756,V253C756,V662C756,V899C756,V1908C756,V2004C756,C756V191,C756V253,C756V662,C756V899,C756V1908,C756V2004,end_cn756);
C757:CNPU6_6 port map (start_cn,clk,rst,V192C757,V254C757,V663C757,V900C757,V1909C757,V2005C757,C757V192,C757V254,C757V663,C757V900,C757V1909,C757V2005,end_cn757);
C758:CNPU6_6 port map (start_cn,clk,rst,V97C758,V255C758,V664C758,V901C758,V1910C758,V2006C758,C758V97,C758V255,C758V664,C758V901,C758V1910,C758V2006,end_cn758);
C759:CNPU6_6 port map (start_cn,clk,rst,V98C759,V256C759,V665C759,V902C759,V1911C759,V2007C759,C759V98,C759V256,C759V665,C759V902,C759V1911,C759V2007,end_cn759);
C760:CNPU6_6 port map (start_cn,clk,rst,V99C760,V257C760,V666C760,V903C760,V1912C760,V2008C760,C760V99,C760V257,C760V666,C760V903,C760V1912,C760V2008,end_cn760);
C761:CNPU6_6 port map (start_cn,clk,rst,V100C761,V258C761,V667C761,V904C761,V1913C761,V2009C761,C761V100,C761V258,C761V667,C761V904,C761V1913,C761V2009,end_cn761);
C762:CNPU6_6 port map (start_cn,clk,rst,V101C762,V259C762,V668C762,V905C762,V1914C762,V2010C762,C762V101,C762V259,C762V668,C762V905,C762V1914,C762V2010,end_cn762);
C763:CNPU6_6 port map (start_cn,clk,rst,V102C763,V260C763,V669C763,V906C763,V1915C763,V2011C763,C763V102,C763V260,C763V669,C763V906,C763V1915,C763V2011,end_cn763);
C764:CNPU6_6 port map (start_cn,clk,rst,V103C764,V261C764,V670C764,V907C764,V1916C764,V2012C764,C764V103,C764V261,C764V670,C764V907,C764V1916,C764V2012,end_cn764);
C765:CNPU6_6 port map (start_cn,clk,rst,V104C765,V262C765,V671C765,V908C765,V1917C765,V2013C765,C765V104,C765V262,C765V671,C765V908,C765V1917,C765V2013,end_cn765);
C766:CNPU6_6 port map (start_cn,clk,rst,V105C766,V263C766,V672C766,V909C766,V1918C766,V2014C766,C766V105,C766V263,C766V672,C766V909,C766V1918,C766V2014,end_cn766);
C767:CNPU6_6 port map (start_cn,clk,rst,V106C767,V264C767,V577C767,V910C767,V1919C767,V2015C767,C767V106,C767V264,C767V577,C767V910,C767V1919,C767V2015,end_cn767);
C768:CNPU6_6 port map (start_cn,clk,rst,V107C768,V265C768,V578C768,V911C768,V1920C768,V2016C768,C768V107,C768V265,C768V578,C768V911,C768V1920,C768V2016,end_cn768);
C769:CNPU7_7 port map (start_cn,clk,rst,V13C769,V468C769,V505C769,V716C769,V1108C769,V1921C769,V2017C769,C769V13,C769V468,C769V505,C769V716,C769V1108,C769V1921,C769V2017,end_cn769);
C770:CNPU7_7 port map (start_cn,clk,rst,V14C770,V469C770,V506C770,V717C770,V1109C770,V1922C770,V2018C770,C770V14,C770V469,C770V506,C770V717,C770V1109,C770V1922,C770V2018,end_cn770);
C771:CNPU7_7 port map (start_cn,clk,rst,V15C771,V470C771,V507C771,V718C771,V1110C771,V1923C771,V2019C771,C771V15,C771V470,C771V507,C771V718,C771V1110,C771V1923,C771V2019,end_cn771);
C772:CNPU7_7 port map (start_cn,clk,rst,V16C772,V471C772,V508C772,V719C772,V1111C772,V1924C772,V2020C772,C772V16,C772V471,C772V508,C772V719,C772V1111,C772V1924,C772V2020,end_cn772);
C773:CNPU7_7 port map (start_cn,clk,rst,V17C773,V472C773,V509C773,V720C773,V1112C773,V1925C773,V2021C773,C773V17,C773V472,C773V509,C773V720,C773V1112,C773V1925,C773V2021,end_cn773);
C774:CNPU7_7 port map (start_cn,clk,rst,V18C774,V473C774,V510C774,V721C774,V1113C774,V1926C774,V2022C774,C774V18,C774V473,C774V510,C774V721,C774V1113,C774V1926,C774V2022,end_cn774);
C775:CNPU7_7 port map (start_cn,clk,rst,V19C775,V474C775,V511C775,V722C775,V1114C775,V1927C775,V2023C775,C775V19,C775V474,C775V511,C775V722,C775V1114,C775V1927,C775V2023,end_cn775);
C776:CNPU7_7 port map (start_cn,clk,rst,V20C776,V475C776,V512C776,V723C776,V1115C776,V1928C776,V2024C776,C776V20,C776V475,C776V512,C776V723,C776V1115,C776V1928,C776V2024,end_cn776);
C777:CNPU7_7 port map (start_cn,clk,rst,V21C777,V476C777,V513C777,V724C777,V1116C777,V1929C777,V2025C777,C777V21,C777V476,C777V513,C777V724,C777V1116,C777V1929,C777V2025,end_cn777);
C778:CNPU7_7 port map (start_cn,clk,rst,V22C778,V477C778,V514C778,V725C778,V1117C778,V1930C778,V2026C778,C778V22,C778V477,C778V514,C778V725,C778V1117,C778V1930,C778V2026,end_cn778);
C779:CNPU7_7 port map (start_cn,clk,rst,V23C779,V478C779,V515C779,V726C779,V1118C779,V1931C779,V2027C779,C779V23,C779V478,C779V515,C779V726,C779V1118,C779V1931,C779V2027,end_cn779);
C780:CNPU7_7 port map (start_cn,clk,rst,V24C780,V479C780,V516C780,V727C780,V1119C780,V1932C780,V2028C780,C780V24,C780V479,C780V516,C780V727,C780V1119,C780V1932,C780V2028,end_cn780);
C781:CNPU7_7 port map (start_cn,clk,rst,V25C781,V480C781,V517C781,V728C781,V1120C781,V1933C781,V2029C781,C781V25,C781V480,C781V517,C781V728,C781V1120,C781V1933,C781V2029,end_cn781);
C782:CNPU7_7 port map (start_cn,clk,rst,V26C782,V385C782,V518C782,V729C782,V1121C782,V1934C782,V2030C782,C782V26,C782V385,C782V518,C782V729,C782V1121,C782V1934,C782V2030,end_cn782);
C783:CNPU7_7 port map (start_cn,clk,rst,V27C783,V386C783,V519C783,V730C783,V1122C783,V1935C783,V2031C783,C783V27,C783V386,C783V519,C783V730,C783V1122,C783V1935,C783V2031,end_cn783);
C784:CNPU7_7 port map (start_cn,clk,rst,V28C784,V387C784,V520C784,V731C784,V1123C784,V1936C784,V2032C784,C784V28,C784V387,C784V520,C784V731,C784V1123,C784V1936,C784V2032,end_cn784);
C785:CNPU7_7 port map (start_cn,clk,rst,V29C785,V388C785,V521C785,V732C785,V1124C785,V1937C785,V2033C785,C785V29,C785V388,C785V521,C785V732,C785V1124,C785V1937,C785V2033,end_cn785);
C786:CNPU7_7 port map (start_cn,clk,rst,V30C786,V389C786,V522C786,V733C786,V1125C786,V1938C786,V2034C786,C786V30,C786V389,C786V522,C786V733,C786V1125,C786V1938,C786V2034,end_cn786);
C787:CNPU7_7 port map (start_cn,clk,rst,V31C787,V390C787,V523C787,V734C787,V1126C787,V1939C787,V2035C787,C787V31,C787V390,C787V523,C787V734,C787V1126,C787V1939,C787V2035,end_cn787);
C788:CNPU7_7 port map (start_cn,clk,rst,V32C788,V391C788,V524C788,V735C788,V1127C788,V1940C788,V2036C788,C788V32,C788V391,C788V524,C788V735,C788V1127,C788V1940,C788V2036,end_cn788);
C789:CNPU7_7 port map (start_cn,clk,rst,V33C789,V392C789,V525C789,V736C789,V1128C789,V1941C789,V2037C789,C789V33,C789V392,C789V525,C789V736,C789V1128,C789V1941,C789V2037,end_cn789);
C790:CNPU7_7 port map (start_cn,clk,rst,V34C790,V393C790,V526C790,V737C790,V1129C790,V1942C790,V2038C790,C790V34,C790V393,C790V526,C790V737,C790V1129,C790V1942,C790V2038,end_cn790);
C791:CNPU7_7 port map (start_cn,clk,rst,V35C791,V394C791,V527C791,V738C791,V1130C791,V1943C791,V2039C791,C791V35,C791V394,C791V527,C791V738,C791V1130,C791V1943,C791V2039,end_cn791);
C792:CNPU7_7 port map (start_cn,clk,rst,V36C792,V395C792,V528C792,V739C792,V1131C792,V1944C792,V2040C792,C792V36,C792V395,C792V528,C792V739,C792V1131,C792V1944,C792V2040,end_cn792);
C793:CNPU7_7 port map (start_cn,clk,rst,V37C793,V396C793,V529C793,V740C793,V1132C793,V1945C793,V2041C793,C793V37,C793V396,C793V529,C793V740,C793V1132,C793V1945,C793V2041,end_cn793);
C794:CNPU7_7 port map (start_cn,clk,rst,V38C794,V397C794,V530C794,V741C794,V1133C794,V1946C794,V2042C794,C794V38,C794V397,C794V530,C794V741,C794V1133,C794V1946,C794V2042,end_cn794);
C795:CNPU7_7 port map (start_cn,clk,rst,V39C795,V398C795,V531C795,V742C795,V1134C795,V1947C795,V2043C795,C795V39,C795V398,C795V531,C795V742,C795V1134,C795V1947,C795V2043,end_cn795);
C796:CNPU7_7 port map (start_cn,clk,rst,V40C796,V399C796,V532C796,V743C796,V1135C796,V1948C796,V2044C796,C796V40,C796V399,C796V532,C796V743,C796V1135,C796V1948,C796V2044,end_cn796);
C797:CNPU7_7 port map (start_cn,clk,rst,V41C797,V400C797,V533C797,V744C797,V1136C797,V1949C797,V2045C797,C797V41,C797V400,C797V533,C797V744,C797V1136,C797V1949,C797V2045,end_cn797);
C798:CNPU7_7 port map (start_cn,clk,rst,V42C798,V401C798,V534C798,V745C798,V1137C798,V1950C798,V2046C798,C798V42,C798V401,C798V534,C798V745,C798V1137,C798V1950,C798V2046,end_cn798);
C799:CNPU7_7 port map (start_cn,clk,rst,V43C799,V402C799,V535C799,V746C799,V1138C799,V1951C799,V2047C799,C799V43,C799V402,C799V535,C799V746,C799V1138,C799V1951,C799V2047,end_cn799);
C800:CNPU7_7 port map (start_cn,clk,rst,V44C800,V403C800,V536C800,V747C800,V1139C800,V1952C800,V2048C800,C800V44,C800V403,C800V536,C800V747,C800V1139,C800V1952,C800V2048,end_cn800);
C801:CNPU7_7 port map (start_cn,clk,rst,V45C801,V404C801,V537C801,V748C801,V1140C801,V1953C801,V2049C801,C801V45,C801V404,C801V537,C801V748,C801V1140,C801V1953,C801V2049,end_cn801);
C802:CNPU7_7 port map (start_cn,clk,rst,V46C802,V405C802,V538C802,V749C802,V1141C802,V1954C802,V2050C802,C802V46,C802V405,C802V538,C802V749,C802V1141,C802V1954,C802V2050,end_cn802);
C803:CNPU7_7 port map (start_cn,clk,rst,V47C803,V406C803,V539C803,V750C803,V1142C803,V1955C803,V2051C803,C803V47,C803V406,C803V539,C803V750,C803V1142,C803V1955,C803V2051,end_cn803);
C804:CNPU7_7 port map (start_cn,clk,rst,V48C804,V407C804,V540C804,V751C804,V1143C804,V1956C804,V2052C804,C804V48,C804V407,C804V540,C804V751,C804V1143,C804V1956,C804V2052,end_cn804);
C805:CNPU7_7 port map (start_cn,clk,rst,V49C805,V408C805,V541C805,V752C805,V1144C805,V1957C805,V2053C805,C805V49,C805V408,C805V541,C805V752,C805V1144,C805V1957,C805V2053,end_cn805);
C806:CNPU7_7 port map (start_cn,clk,rst,V50C806,V409C806,V542C806,V753C806,V1145C806,V1958C806,V2054C806,C806V50,C806V409,C806V542,C806V753,C806V1145,C806V1958,C806V2054,end_cn806);
C807:CNPU7_7 port map (start_cn,clk,rst,V51C807,V410C807,V543C807,V754C807,V1146C807,V1959C807,V2055C807,C807V51,C807V410,C807V543,C807V754,C807V1146,C807V1959,C807V2055,end_cn807);
C808:CNPU7_7 port map (start_cn,clk,rst,V52C808,V411C808,V544C808,V755C808,V1147C808,V1960C808,V2056C808,C808V52,C808V411,C808V544,C808V755,C808V1147,C808V1960,C808V2056,end_cn808);
C809:CNPU7_7 port map (start_cn,clk,rst,V53C809,V412C809,V545C809,V756C809,V1148C809,V1961C809,V2057C809,C809V53,C809V412,C809V545,C809V756,C809V1148,C809V1961,C809V2057,end_cn809);
C810:CNPU7_7 port map (start_cn,clk,rst,V54C810,V413C810,V546C810,V757C810,V1149C810,V1962C810,V2058C810,C810V54,C810V413,C810V546,C810V757,C810V1149,C810V1962,C810V2058,end_cn810);
C811:CNPU7_7 port map (start_cn,clk,rst,V55C811,V414C811,V547C811,V758C811,V1150C811,V1963C811,V2059C811,C811V55,C811V414,C811V547,C811V758,C811V1150,C811V1963,C811V2059,end_cn811);
C812:CNPU7_7 port map (start_cn,clk,rst,V56C812,V415C812,V548C812,V759C812,V1151C812,V1964C812,V2060C812,C812V56,C812V415,C812V548,C812V759,C812V1151,C812V1964,C812V2060,end_cn812);
C813:CNPU7_7 port map (start_cn,clk,rst,V57C813,V416C813,V549C813,V760C813,V1152C813,V1965C813,V2061C813,C813V57,C813V416,C813V549,C813V760,C813V1152,C813V1965,C813V2061,end_cn813);
C814:CNPU7_7 port map (start_cn,clk,rst,V58C814,V417C814,V550C814,V761C814,V1057C814,V1966C814,V2062C814,C814V58,C814V417,C814V550,C814V761,C814V1057,C814V1966,C814V2062,end_cn814);
C815:CNPU7_7 port map (start_cn,clk,rst,V59C815,V418C815,V551C815,V762C815,V1058C815,V1967C815,V2063C815,C815V59,C815V418,C815V551,C815V762,C815V1058,C815V1967,C815V2063,end_cn815);
C816:CNPU7_7 port map (start_cn,clk,rst,V60C816,V419C816,V552C816,V763C816,V1059C816,V1968C816,V2064C816,C816V60,C816V419,C816V552,C816V763,C816V1059,C816V1968,C816V2064,end_cn816);
C817:CNPU7_7 port map (start_cn,clk,rst,V61C817,V420C817,V553C817,V764C817,V1060C817,V1969C817,V2065C817,C817V61,C817V420,C817V553,C817V764,C817V1060,C817V1969,C817V2065,end_cn817);
C818:CNPU7_7 port map (start_cn,clk,rst,V62C818,V421C818,V554C818,V765C818,V1061C818,V1970C818,V2066C818,C818V62,C818V421,C818V554,C818V765,C818V1061,C818V1970,C818V2066,end_cn818);
C819:CNPU7_7 port map (start_cn,clk,rst,V63C819,V422C819,V555C819,V766C819,V1062C819,V1971C819,V2067C819,C819V63,C819V422,C819V555,C819V766,C819V1062,C819V1971,C819V2067,end_cn819);
C820:CNPU7_7 port map (start_cn,clk,rst,V64C820,V423C820,V556C820,V767C820,V1063C820,V1972C820,V2068C820,C820V64,C820V423,C820V556,C820V767,C820V1063,C820V1972,C820V2068,end_cn820);
C821:CNPU7_7 port map (start_cn,clk,rst,V65C821,V424C821,V557C821,V768C821,V1064C821,V1973C821,V2069C821,C821V65,C821V424,C821V557,C821V768,C821V1064,C821V1973,C821V2069,end_cn821);
C822:CNPU7_7 port map (start_cn,clk,rst,V66C822,V425C822,V558C822,V673C822,V1065C822,V1974C822,V2070C822,C822V66,C822V425,C822V558,C822V673,C822V1065,C822V1974,C822V2070,end_cn822);
C823:CNPU7_7 port map (start_cn,clk,rst,V67C823,V426C823,V559C823,V674C823,V1066C823,V1975C823,V2071C823,C823V67,C823V426,C823V559,C823V674,C823V1066,C823V1975,C823V2071,end_cn823);
C824:CNPU7_7 port map (start_cn,clk,rst,V68C824,V427C824,V560C824,V675C824,V1067C824,V1976C824,V2072C824,C824V68,C824V427,C824V560,C824V675,C824V1067,C824V1976,C824V2072,end_cn824);
C825:CNPU7_7 port map (start_cn,clk,rst,V69C825,V428C825,V561C825,V676C825,V1068C825,V1977C825,V2073C825,C825V69,C825V428,C825V561,C825V676,C825V1068,C825V1977,C825V2073,end_cn825);
C826:CNPU7_7 port map (start_cn,clk,rst,V70C826,V429C826,V562C826,V677C826,V1069C826,V1978C826,V2074C826,C826V70,C826V429,C826V562,C826V677,C826V1069,C826V1978,C826V2074,end_cn826);
C827:CNPU7_7 port map (start_cn,clk,rst,V71C827,V430C827,V563C827,V678C827,V1070C827,V1979C827,V2075C827,C827V71,C827V430,C827V563,C827V678,C827V1070,C827V1979,C827V2075,end_cn827);
C828:CNPU7_7 port map (start_cn,clk,rst,V72C828,V431C828,V564C828,V679C828,V1071C828,V1980C828,V2076C828,C828V72,C828V431,C828V564,C828V679,C828V1071,C828V1980,C828V2076,end_cn828);
C829:CNPU7_7 port map (start_cn,clk,rst,V73C829,V432C829,V565C829,V680C829,V1072C829,V1981C829,V2077C829,C829V73,C829V432,C829V565,C829V680,C829V1072,C829V1981,C829V2077,end_cn829);
C830:CNPU7_7 port map (start_cn,clk,rst,V74C830,V433C830,V566C830,V681C830,V1073C830,V1982C830,V2078C830,C830V74,C830V433,C830V566,C830V681,C830V1073,C830V1982,C830V2078,end_cn830);
C831:CNPU7_7 port map (start_cn,clk,rst,V75C831,V434C831,V567C831,V682C831,V1074C831,V1983C831,V2079C831,C831V75,C831V434,C831V567,C831V682,C831V1074,C831V1983,C831V2079,end_cn831);
C832:CNPU7_7 port map (start_cn,clk,rst,V76C832,V435C832,V568C832,V683C832,V1075C832,V1984C832,V2080C832,C832V76,C832V435,C832V568,C832V683,C832V1075,C832V1984,C832V2080,end_cn832);
C833:CNPU7_7 port map (start_cn,clk,rst,V77C833,V436C833,V569C833,V684C833,V1076C833,V1985C833,V2081C833,C833V77,C833V436,C833V569,C833V684,C833V1076,C833V1985,C833V2081,end_cn833);
C834:CNPU7_7 port map (start_cn,clk,rst,V78C834,V437C834,V570C834,V685C834,V1077C834,V1986C834,V2082C834,C834V78,C834V437,C834V570,C834V685,C834V1077,C834V1986,C834V2082,end_cn834);
C835:CNPU7_7 port map (start_cn,clk,rst,V79C835,V438C835,V571C835,V686C835,V1078C835,V1987C835,V2083C835,C835V79,C835V438,C835V571,C835V686,C835V1078,C835V1987,C835V2083,end_cn835);
C836:CNPU7_7 port map (start_cn,clk,rst,V80C836,V439C836,V572C836,V687C836,V1079C836,V1988C836,V2084C836,C836V80,C836V439,C836V572,C836V687,C836V1079,C836V1988,C836V2084,end_cn836);
C837:CNPU7_7 port map (start_cn,clk,rst,V81C837,V440C837,V573C837,V688C837,V1080C837,V1989C837,V2085C837,C837V81,C837V440,C837V573,C837V688,C837V1080,C837V1989,C837V2085,end_cn837);
C838:CNPU7_7 port map (start_cn,clk,rst,V82C838,V441C838,V574C838,V689C838,V1081C838,V1990C838,V2086C838,C838V82,C838V441,C838V574,C838V689,C838V1081,C838V1990,C838V2086,end_cn838);
C839:CNPU7_7 port map (start_cn,clk,rst,V83C839,V442C839,V575C839,V690C839,V1082C839,V1991C839,V2087C839,C839V83,C839V442,C839V575,C839V690,C839V1082,C839V1991,C839V2087,end_cn839);
C840:CNPU7_7 port map (start_cn,clk,rst,V84C840,V443C840,V576C840,V691C840,V1083C840,V1992C840,V2088C840,C840V84,C840V443,C840V576,C840V691,C840V1083,C840V1992,C840V2088,end_cn840);
C841:CNPU7_7 port map (start_cn,clk,rst,V85C841,V444C841,V481C841,V692C841,V1084C841,V1993C841,V2089C841,C841V85,C841V444,C841V481,C841V692,C841V1084,C841V1993,C841V2089,end_cn841);
C842:CNPU7_7 port map (start_cn,clk,rst,V86C842,V445C842,V482C842,V693C842,V1085C842,V1994C842,V2090C842,C842V86,C842V445,C842V482,C842V693,C842V1085,C842V1994,C842V2090,end_cn842);
C843:CNPU7_7 port map (start_cn,clk,rst,V87C843,V446C843,V483C843,V694C843,V1086C843,V1995C843,V2091C843,C843V87,C843V446,C843V483,C843V694,C843V1086,C843V1995,C843V2091,end_cn843);
C844:CNPU7_7 port map (start_cn,clk,rst,V88C844,V447C844,V484C844,V695C844,V1087C844,V1996C844,V2092C844,C844V88,C844V447,C844V484,C844V695,C844V1087,C844V1996,C844V2092,end_cn844);
C845:CNPU7_7 port map (start_cn,clk,rst,V89C845,V448C845,V485C845,V696C845,V1088C845,V1997C845,V2093C845,C845V89,C845V448,C845V485,C845V696,C845V1088,C845V1997,C845V2093,end_cn845);
C846:CNPU7_7 port map (start_cn,clk,rst,V90C846,V449C846,V486C846,V697C846,V1089C846,V1998C846,V2094C846,C846V90,C846V449,C846V486,C846V697,C846V1089,C846V1998,C846V2094,end_cn846);
C847:CNPU7_7 port map (start_cn,clk,rst,V91C847,V450C847,V487C847,V698C847,V1090C847,V1999C847,V2095C847,C847V91,C847V450,C847V487,C847V698,C847V1090,C847V1999,C847V2095,end_cn847);
C848:CNPU7_7 port map (start_cn,clk,rst,V92C848,V451C848,V488C848,V699C848,V1091C848,V2000C848,V2096C848,C848V92,C848V451,C848V488,C848V699,C848V1091,C848V2000,C848V2096,end_cn848);
C849:CNPU7_7 port map (start_cn,clk,rst,V93C849,V452C849,V489C849,V700C849,V1092C849,V2001C849,V2097C849,C849V93,C849V452,C849V489,C849V700,C849V1092,C849V2001,C849V2097,end_cn849);
C850:CNPU7_7 port map (start_cn,clk,rst,V94C850,V453C850,V490C850,V701C850,V1093C850,V2002C850,V2098C850,C850V94,C850V453,C850V490,C850V701,C850V1093,C850V2002,C850V2098,end_cn850);
C851:CNPU7_7 port map (start_cn,clk,rst,V95C851,V454C851,V491C851,V702C851,V1094C851,V2003C851,V2099C851,C851V95,C851V454,C851V491,C851V702,C851V1094,C851V2003,C851V2099,end_cn851);
C852:CNPU7_7 port map (start_cn,clk,rst,V96C852,V455C852,V492C852,V703C852,V1095C852,V2004C852,V2100C852,C852V96,C852V455,C852V492,C852V703,C852V1095,C852V2004,C852V2100,end_cn852);
C853:CNPU7_7 port map (start_cn,clk,rst,V1C853,V456C853,V493C853,V704C853,V1096C853,V2005C853,V2101C853,C853V1,C853V456,C853V493,C853V704,C853V1096,C853V2005,C853V2101,end_cn853);
C854:CNPU7_7 port map (start_cn,clk,rst,V2C854,V457C854,V494C854,V705C854,V1097C854,V2006C854,V2102C854,C854V2,C854V457,C854V494,C854V705,C854V1097,C854V2006,C854V2102,end_cn854);
C855:CNPU7_7 port map (start_cn,clk,rst,V3C855,V458C855,V495C855,V706C855,V1098C855,V2007C855,V2103C855,C855V3,C855V458,C855V495,C855V706,C855V1098,C855V2007,C855V2103,end_cn855);
C856:CNPU7_7 port map (start_cn,clk,rst,V4C856,V459C856,V496C856,V707C856,V1099C856,V2008C856,V2104C856,C856V4,C856V459,C856V496,C856V707,C856V1099,C856V2008,C856V2104,end_cn856);
C857:CNPU7_7 port map (start_cn,clk,rst,V5C857,V460C857,V497C857,V708C857,V1100C857,V2009C857,V2105C857,C857V5,C857V460,C857V497,C857V708,C857V1100,C857V2009,C857V2105,end_cn857);
C858:CNPU7_7 port map (start_cn,clk,rst,V6C858,V461C858,V498C858,V709C858,V1101C858,V2010C858,V2106C858,C858V6,C858V461,C858V498,C858V709,C858V1101,C858V2010,C858V2106,end_cn858);
C859:CNPU7_7 port map (start_cn,clk,rst,V7C859,V462C859,V499C859,V710C859,V1102C859,V2011C859,V2107C859,C859V7,C859V462,C859V499,C859V710,C859V1102,C859V2011,C859V2107,end_cn859);
C860:CNPU7_7 port map (start_cn,clk,rst,V8C860,V463C860,V500C860,V711C860,V1103C860,V2012C860,V2108C860,C860V8,C860V463,C860V500,C860V711,C860V1103,C860V2012,C860V2108,end_cn860);
C861:CNPU7_7 port map (start_cn,clk,rst,V9C861,V464C861,V501C861,V712C861,V1104C861,V2013C861,V2109C861,C861V9,C861V464,C861V501,C861V712,C861V1104,C861V2013,C861V2109,end_cn861);
C862:CNPU7_7 port map (start_cn,clk,rst,V10C862,V465C862,V502C862,V713C862,V1105C862,V2014C862,V2110C862,C862V10,C862V465,C862V502,C862V713,C862V1105,C862V2014,C862V2110,end_cn862);
C863:CNPU7_7 port map (start_cn,clk,rst,V11C863,V466C863,V503C863,V714C863,V1106C863,V2015C863,V2111C863,C863V11,C863V466,C863V503,C863V714,C863V1106,C863V2015,C863V2111,end_cn863);
C864:CNPU7_7 port map (start_cn,clk,rst,V12C864,V467C864,V504C864,V715C864,V1107C864,V2016C864,V2112C864,C864V12,C864V467,C864V504,C864V715,C864V1107,C864V2016,C864V2112,end_cn864);
C865:CNPU6_6 port map (start_cn,clk,rst,V575C865,V732C865,V1031C865,V1129C865,V2017C865,V2113C865,C865V575,C865V732,C865V1031,C865V1129,C865V2017,C865V2113,end_cn865);
C866:CNPU6_6 port map (start_cn,clk,rst,V576C866,V733C866,V1032C866,V1130C866,V2018C866,V2114C866,C866V576,C866V733,C866V1032,C866V1130,C866V2018,C866V2114,end_cn866);
C867:CNPU6_6 port map (start_cn,clk,rst,V481C867,V734C867,V1033C867,V1131C867,V2019C867,V2115C867,C867V481,C867V734,C867V1033,C867V1131,C867V2019,C867V2115,end_cn867);
C868:CNPU6_6 port map (start_cn,clk,rst,V482C868,V735C868,V1034C868,V1132C868,V2020C868,V2116C868,C868V482,C868V735,C868V1034,C868V1132,C868V2020,C868V2116,end_cn868);
C869:CNPU6_6 port map (start_cn,clk,rst,V483C869,V736C869,V1035C869,V1133C869,V2021C869,V2117C869,C869V483,C869V736,C869V1035,C869V1133,C869V2021,C869V2117,end_cn869);
C870:CNPU6_6 port map (start_cn,clk,rst,V484C870,V737C870,V1036C870,V1134C870,V2022C870,V2118C870,C870V484,C870V737,C870V1036,C870V1134,C870V2022,C870V2118,end_cn870);
C871:CNPU6_6 port map (start_cn,clk,rst,V485C871,V738C871,V1037C871,V1135C871,V2023C871,V2119C871,C871V485,C871V738,C871V1037,C871V1135,C871V2023,C871V2119,end_cn871);
C872:CNPU6_6 port map (start_cn,clk,rst,V486C872,V739C872,V1038C872,V1136C872,V2024C872,V2120C872,C872V486,C872V739,C872V1038,C872V1136,C872V2024,C872V2120,end_cn872);
C873:CNPU6_6 port map (start_cn,clk,rst,V487C873,V740C873,V1039C873,V1137C873,V2025C873,V2121C873,C873V487,C873V740,C873V1039,C873V1137,C873V2025,C873V2121,end_cn873);
C874:CNPU6_6 port map (start_cn,clk,rst,V488C874,V741C874,V1040C874,V1138C874,V2026C874,V2122C874,C874V488,C874V741,C874V1040,C874V1138,C874V2026,C874V2122,end_cn874);
C875:CNPU6_6 port map (start_cn,clk,rst,V489C875,V742C875,V1041C875,V1139C875,V2027C875,V2123C875,C875V489,C875V742,C875V1041,C875V1139,C875V2027,C875V2123,end_cn875);
C876:CNPU6_6 port map (start_cn,clk,rst,V490C876,V743C876,V1042C876,V1140C876,V2028C876,V2124C876,C876V490,C876V743,C876V1042,C876V1140,C876V2028,C876V2124,end_cn876);
C877:CNPU6_6 port map (start_cn,clk,rst,V491C877,V744C877,V1043C877,V1141C877,V2029C877,V2125C877,C877V491,C877V744,C877V1043,C877V1141,C877V2029,C877V2125,end_cn877);
C878:CNPU6_6 port map (start_cn,clk,rst,V492C878,V745C878,V1044C878,V1142C878,V2030C878,V2126C878,C878V492,C878V745,C878V1044,C878V1142,C878V2030,C878V2126,end_cn878);
C879:CNPU6_6 port map (start_cn,clk,rst,V493C879,V746C879,V1045C879,V1143C879,V2031C879,V2127C879,C879V493,C879V746,C879V1045,C879V1143,C879V2031,C879V2127,end_cn879);
C880:CNPU6_6 port map (start_cn,clk,rst,V494C880,V747C880,V1046C880,V1144C880,V2032C880,V2128C880,C880V494,C880V747,C880V1046,C880V1144,C880V2032,C880V2128,end_cn880);
C881:CNPU6_6 port map (start_cn,clk,rst,V495C881,V748C881,V1047C881,V1145C881,V2033C881,V2129C881,C881V495,C881V748,C881V1047,C881V1145,C881V2033,C881V2129,end_cn881);
C882:CNPU6_6 port map (start_cn,clk,rst,V496C882,V749C882,V1048C882,V1146C882,V2034C882,V2130C882,C882V496,C882V749,C882V1048,C882V1146,C882V2034,C882V2130,end_cn882);
C883:CNPU6_6 port map (start_cn,clk,rst,V497C883,V750C883,V1049C883,V1147C883,V2035C883,V2131C883,C883V497,C883V750,C883V1049,C883V1147,C883V2035,C883V2131,end_cn883);
C884:CNPU6_6 port map (start_cn,clk,rst,V498C884,V751C884,V1050C884,V1148C884,V2036C884,V2132C884,C884V498,C884V751,C884V1050,C884V1148,C884V2036,C884V2132,end_cn884);
C885:CNPU6_6 port map (start_cn,clk,rst,V499C885,V752C885,V1051C885,V1149C885,V2037C885,V2133C885,C885V499,C885V752,C885V1051,C885V1149,C885V2037,C885V2133,end_cn885);
C886:CNPU6_6 port map (start_cn,clk,rst,V500C886,V753C886,V1052C886,V1150C886,V2038C886,V2134C886,C886V500,C886V753,C886V1052,C886V1150,C886V2038,C886V2134,end_cn886);
C887:CNPU6_6 port map (start_cn,clk,rst,V501C887,V754C887,V1053C887,V1151C887,V2039C887,V2135C887,C887V501,C887V754,C887V1053,C887V1151,C887V2039,C887V2135,end_cn887);
C888:CNPU6_6 port map (start_cn,clk,rst,V502C888,V755C888,V1054C888,V1152C888,V2040C888,V2136C888,C888V502,C888V755,C888V1054,C888V1152,C888V2040,C888V2136,end_cn888);
C889:CNPU6_6 port map (start_cn,clk,rst,V503C889,V756C889,V1055C889,V1057C889,V2041C889,V2137C889,C889V503,C889V756,C889V1055,C889V1057,C889V2041,C889V2137,end_cn889);
C890:CNPU6_6 port map (start_cn,clk,rst,V504C890,V757C890,V1056C890,V1058C890,V2042C890,V2138C890,C890V504,C890V757,C890V1056,C890V1058,C890V2042,C890V2138,end_cn890);
C891:CNPU6_6 port map (start_cn,clk,rst,V505C891,V758C891,V961C891,V1059C891,V2043C891,V2139C891,C891V505,C891V758,C891V961,C891V1059,C891V2043,C891V2139,end_cn891);
C892:CNPU6_6 port map (start_cn,clk,rst,V506C892,V759C892,V962C892,V1060C892,V2044C892,V2140C892,C892V506,C892V759,C892V962,C892V1060,C892V2044,C892V2140,end_cn892);
C893:CNPU6_6 port map (start_cn,clk,rst,V507C893,V760C893,V963C893,V1061C893,V2045C893,V2141C893,C893V507,C893V760,C893V963,C893V1061,C893V2045,C893V2141,end_cn893);
C894:CNPU6_6 port map (start_cn,clk,rst,V508C894,V761C894,V964C894,V1062C894,V2046C894,V2142C894,C894V508,C894V761,C894V964,C894V1062,C894V2046,C894V2142,end_cn894);
C895:CNPU6_6 port map (start_cn,clk,rst,V509C895,V762C895,V965C895,V1063C895,V2047C895,V2143C895,C895V509,C895V762,C895V965,C895V1063,C895V2047,C895V2143,end_cn895);
C896:CNPU6_6 port map (start_cn,clk,rst,V510C896,V763C896,V966C896,V1064C896,V2048C896,V2144C896,C896V510,C896V763,C896V966,C896V1064,C896V2048,C896V2144,end_cn896);
C897:CNPU6_6 port map (start_cn,clk,rst,V511C897,V764C897,V967C897,V1065C897,V2049C897,V2145C897,C897V511,C897V764,C897V967,C897V1065,C897V2049,C897V2145,end_cn897);
C898:CNPU6_6 port map (start_cn,clk,rst,V512C898,V765C898,V968C898,V1066C898,V2050C898,V2146C898,C898V512,C898V765,C898V968,C898V1066,C898V2050,C898V2146,end_cn898);
C899:CNPU6_6 port map (start_cn,clk,rst,V513C899,V766C899,V969C899,V1067C899,V2051C899,V2147C899,C899V513,C899V766,C899V969,C899V1067,C899V2051,C899V2147,end_cn899);
C900:CNPU6_6 port map (start_cn,clk,rst,V514C900,V767C900,V970C900,V1068C900,V2052C900,V2148C900,C900V514,C900V767,C900V970,C900V1068,C900V2052,C900V2148,end_cn900);
C901:CNPU6_6 port map (start_cn,clk,rst,V515C901,V768C901,V971C901,V1069C901,V2053C901,V2149C901,C901V515,C901V768,C901V971,C901V1069,C901V2053,C901V2149,end_cn901);
C902:CNPU6_6 port map (start_cn,clk,rst,V516C902,V673C902,V972C902,V1070C902,V2054C902,V2150C902,C902V516,C902V673,C902V972,C902V1070,C902V2054,C902V2150,end_cn902);
C903:CNPU6_6 port map (start_cn,clk,rst,V517C903,V674C903,V973C903,V1071C903,V2055C903,V2151C903,C903V517,C903V674,C903V973,C903V1071,C903V2055,C903V2151,end_cn903);
C904:CNPU6_6 port map (start_cn,clk,rst,V518C904,V675C904,V974C904,V1072C904,V2056C904,V2152C904,C904V518,C904V675,C904V974,C904V1072,C904V2056,C904V2152,end_cn904);
C905:CNPU6_6 port map (start_cn,clk,rst,V519C905,V676C905,V975C905,V1073C905,V2057C905,V2153C905,C905V519,C905V676,C905V975,C905V1073,C905V2057,C905V2153,end_cn905);
C906:CNPU6_6 port map (start_cn,clk,rst,V520C906,V677C906,V976C906,V1074C906,V2058C906,V2154C906,C906V520,C906V677,C906V976,C906V1074,C906V2058,C906V2154,end_cn906);
C907:CNPU6_6 port map (start_cn,clk,rst,V521C907,V678C907,V977C907,V1075C907,V2059C907,V2155C907,C907V521,C907V678,C907V977,C907V1075,C907V2059,C907V2155,end_cn907);
C908:CNPU6_6 port map (start_cn,clk,rst,V522C908,V679C908,V978C908,V1076C908,V2060C908,V2156C908,C908V522,C908V679,C908V978,C908V1076,C908V2060,C908V2156,end_cn908);
C909:CNPU6_6 port map (start_cn,clk,rst,V523C909,V680C909,V979C909,V1077C909,V2061C909,V2157C909,C909V523,C909V680,C909V979,C909V1077,C909V2061,C909V2157,end_cn909);
C910:CNPU6_6 port map (start_cn,clk,rst,V524C910,V681C910,V980C910,V1078C910,V2062C910,V2158C910,C910V524,C910V681,C910V980,C910V1078,C910V2062,C910V2158,end_cn910);
C911:CNPU6_6 port map (start_cn,clk,rst,V525C911,V682C911,V981C911,V1079C911,V2063C911,V2159C911,C911V525,C911V682,C911V981,C911V1079,C911V2063,C911V2159,end_cn911);
C912:CNPU6_6 port map (start_cn,clk,rst,V526C912,V683C912,V982C912,V1080C912,V2064C912,V2160C912,C912V526,C912V683,C912V982,C912V1080,C912V2064,C912V2160,end_cn912);
C913:CNPU6_6 port map (start_cn,clk,rst,V527C913,V684C913,V983C913,V1081C913,V2065C913,V2161C913,C913V527,C913V684,C913V983,C913V1081,C913V2065,C913V2161,end_cn913);
C914:CNPU6_6 port map (start_cn,clk,rst,V528C914,V685C914,V984C914,V1082C914,V2066C914,V2162C914,C914V528,C914V685,C914V984,C914V1082,C914V2066,C914V2162,end_cn914);
C915:CNPU6_6 port map (start_cn,clk,rst,V529C915,V686C915,V985C915,V1083C915,V2067C915,V2163C915,C915V529,C915V686,C915V985,C915V1083,C915V2067,C915V2163,end_cn915);
C916:CNPU6_6 port map (start_cn,clk,rst,V530C916,V687C916,V986C916,V1084C916,V2068C916,V2164C916,C916V530,C916V687,C916V986,C916V1084,C916V2068,C916V2164,end_cn916);
C917:CNPU6_6 port map (start_cn,clk,rst,V531C917,V688C917,V987C917,V1085C917,V2069C917,V2165C917,C917V531,C917V688,C917V987,C917V1085,C917V2069,C917V2165,end_cn917);
C918:CNPU6_6 port map (start_cn,clk,rst,V532C918,V689C918,V988C918,V1086C918,V2070C918,V2166C918,C918V532,C918V689,C918V988,C918V1086,C918V2070,C918V2166,end_cn918);
C919:CNPU6_6 port map (start_cn,clk,rst,V533C919,V690C919,V989C919,V1087C919,V2071C919,V2167C919,C919V533,C919V690,C919V989,C919V1087,C919V2071,C919V2167,end_cn919);
C920:CNPU6_6 port map (start_cn,clk,rst,V534C920,V691C920,V990C920,V1088C920,V2072C920,V2168C920,C920V534,C920V691,C920V990,C920V1088,C920V2072,C920V2168,end_cn920);
C921:CNPU6_6 port map (start_cn,clk,rst,V535C921,V692C921,V991C921,V1089C921,V2073C921,V2169C921,C921V535,C921V692,C921V991,C921V1089,C921V2073,C921V2169,end_cn921);
C922:CNPU6_6 port map (start_cn,clk,rst,V536C922,V693C922,V992C922,V1090C922,V2074C922,V2170C922,C922V536,C922V693,C922V992,C922V1090,C922V2074,C922V2170,end_cn922);
C923:CNPU6_6 port map (start_cn,clk,rst,V537C923,V694C923,V993C923,V1091C923,V2075C923,V2171C923,C923V537,C923V694,C923V993,C923V1091,C923V2075,C923V2171,end_cn923);
C924:CNPU6_6 port map (start_cn,clk,rst,V538C924,V695C924,V994C924,V1092C924,V2076C924,V2172C924,C924V538,C924V695,C924V994,C924V1092,C924V2076,C924V2172,end_cn924);
C925:CNPU6_6 port map (start_cn,clk,rst,V539C925,V696C925,V995C925,V1093C925,V2077C925,V2173C925,C925V539,C925V696,C925V995,C925V1093,C925V2077,C925V2173,end_cn925);
C926:CNPU6_6 port map (start_cn,clk,rst,V540C926,V697C926,V996C926,V1094C926,V2078C926,V2174C926,C926V540,C926V697,C926V996,C926V1094,C926V2078,C926V2174,end_cn926);
C927:CNPU6_6 port map (start_cn,clk,rst,V541C927,V698C927,V997C927,V1095C927,V2079C927,V2175C927,C927V541,C927V698,C927V997,C927V1095,C927V2079,C927V2175,end_cn927);
C928:CNPU6_6 port map (start_cn,clk,rst,V542C928,V699C928,V998C928,V1096C928,V2080C928,V2176C928,C928V542,C928V699,C928V998,C928V1096,C928V2080,C928V2176,end_cn928);
C929:CNPU6_6 port map (start_cn,clk,rst,V543C929,V700C929,V999C929,V1097C929,V2081C929,V2177C929,C929V543,C929V700,C929V999,C929V1097,C929V2081,C929V2177,end_cn929);
C930:CNPU6_6 port map (start_cn,clk,rst,V544C930,V701C930,V1000C930,V1098C930,V2082C930,V2178C930,C930V544,C930V701,C930V1000,C930V1098,C930V2082,C930V2178,end_cn930);
C931:CNPU6_6 port map (start_cn,clk,rst,V545C931,V702C931,V1001C931,V1099C931,V2083C931,V2179C931,C931V545,C931V702,C931V1001,C931V1099,C931V2083,C931V2179,end_cn931);
C932:CNPU6_6 port map (start_cn,clk,rst,V546C932,V703C932,V1002C932,V1100C932,V2084C932,V2180C932,C932V546,C932V703,C932V1002,C932V1100,C932V2084,C932V2180,end_cn932);
C933:CNPU6_6 port map (start_cn,clk,rst,V547C933,V704C933,V1003C933,V1101C933,V2085C933,V2181C933,C933V547,C933V704,C933V1003,C933V1101,C933V2085,C933V2181,end_cn933);
C934:CNPU6_6 port map (start_cn,clk,rst,V548C934,V705C934,V1004C934,V1102C934,V2086C934,V2182C934,C934V548,C934V705,C934V1004,C934V1102,C934V2086,C934V2182,end_cn934);
C935:CNPU6_6 port map (start_cn,clk,rst,V549C935,V706C935,V1005C935,V1103C935,V2087C935,V2183C935,C935V549,C935V706,C935V1005,C935V1103,C935V2087,C935V2183,end_cn935);
C936:CNPU6_6 port map (start_cn,clk,rst,V550C936,V707C936,V1006C936,V1104C936,V2088C936,V2184C936,C936V550,C936V707,C936V1006,C936V1104,C936V2088,C936V2184,end_cn936);
C937:CNPU6_6 port map (start_cn,clk,rst,V551C937,V708C937,V1007C937,V1105C937,V2089C937,V2185C937,C937V551,C937V708,C937V1007,C937V1105,C937V2089,C937V2185,end_cn937);
C938:CNPU6_6 port map (start_cn,clk,rst,V552C938,V709C938,V1008C938,V1106C938,V2090C938,V2186C938,C938V552,C938V709,C938V1008,C938V1106,C938V2090,C938V2186,end_cn938);
C939:CNPU6_6 port map (start_cn,clk,rst,V553C939,V710C939,V1009C939,V1107C939,V2091C939,V2187C939,C939V553,C939V710,C939V1009,C939V1107,C939V2091,C939V2187,end_cn939);
C940:CNPU6_6 port map (start_cn,clk,rst,V554C940,V711C940,V1010C940,V1108C940,V2092C940,V2188C940,C940V554,C940V711,C940V1010,C940V1108,C940V2092,C940V2188,end_cn940);
C941:CNPU6_6 port map (start_cn,clk,rst,V555C941,V712C941,V1011C941,V1109C941,V2093C941,V2189C941,C941V555,C941V712,C941V1011,C941V1109,C941V2093,C941V2189,end_cn941);
C942:CNPU6_6 port map (start_cn,clk,rst,V556C942,V713C942,V1012C942,V1110C942,V2094C942,V2190C942,C942V556,C942V713,C942V1012,C942V1110,C942V2094,C942V2190,end_cn942);
C943:CNPU6_6 port map (start_cn,clk,rst,V557C943,V714C943,V1013C943,V1111C943,V2095C943,V2191C943,C943V557,C943V714,C943V1013,C943V1111,C943V2095,C943V2191,end_cn943);
C944:CNPU6_6 port map (start_cn,clk,rst,V558C944,V715C944,V1014C944,V1112C944,V2096C944,V2192C944,C944V558,C944V715,C944V1014,C944V1112,C944V2096,C944V2192,end_cn944);
C945:CNPU6_6 port map (start_cn,clk,rst,V559C945,V716C945,V1015C945,V1113C945,V2097C945,V2193C945,C945V559,C945V716,C945V1015,C945V1113,C945V2097,C945V2193,end_cn945);
C946:CNPU6_6 port map (start_cn,clk,rst,V560C946,V717C946,V1016C946,V1114C946,V2098C946,V2194C946,C946V560,C946V717,C946V1016,C946V1114,C946V2098,C946V2194,end_cn946);
C947:CNPU6_6 port map (start_cn,clk,rst,V561C947,V718C947,V1017C947,V1115C947,V2099C947,V2195C947,C947V561,C947V718,C947V1017,C947V1115,C947V2099,C947V2195,end_cn947);
C948:CNPU6_6 port map (start_cn,clk,rst,V562C948,V719C948,V1018C948,V1116C948,V2100C948,V2196C948,C948V562,C948V719,C948V1018,C948V1116,C948V2100,C948V2196,end_cn948);
C949:CNPU6_6 port map (start_cn,clk,rst,V563C949,V720C949,V1019C949,V1117C949,V2101C949,V2197C949,C949V563,C949V720,C949V1019,C949V1117,C949V2101,C949V2197,end_cn949);
C950:CNPU6_6 port map (start_cn,clk,rst,V564C950,V721C950,V1020C950,V1118C950,V2102C950,V2198C950,C950V564,C950V721,C950V1020,C950V1118,C950V2102,C950V2198,end_cn950);
C951:CNPU6_6 port map (start_cn,clk,rst,V565C951,V722C951,V1021C951,V1119C951,V2103C951,V2199C951,C951V565,C951V722,C951V1021,C951V1119,C951V2103,C951V2199,end_cn951);
C952:CNPU6_6 port map (start_cn,clk,rst,V566C952,V723C952,V1022C952,V1120C952,V2104C952,V2200C952,C952V566,C952V723,C952V1022,C952V1120,C952V2104,C952V2200,end_cn952);
C953:CNPU6_6 port map (start_cn,clk,rst,V567C953,V724C953,V1023C953,V1121C953,V2105C953,V2201C953,C953V567,C953V724,C953V1023,C953V1121,C953V2105,C953V2201,end_cn953);
C954:CNPU6_6 port map (start_cn,clk,rst,V568C954,V725C954,V1024C954,V1122C954,V2106C954,V2202C954,C954V568,C954V725,C954V1024,C954V1122,C954V2106,C954V2202,end_cn954);
C955:CNPU6_6 port map (start_cn,clk,rst,V569C955,V726C955,V1025C955,V1123C955,V2107C955,V2203C955,C955V569,C955V726,C955V1025,C955V1123,C955V2107,C955V2203,end_cn955);
C956:CNPU6_6 port map (start_cn,clk,rst,V570C956,V727C956,V1026C956,V1124C956,V2108C956,V2204C956,C956V570,C956V727,C956V1026,C956V1124,C956V2108,C956V2204,end_cn956);
C957:CNPU6_6 port map (start_cn,clk,rst,V571C957,V728C957,V1027C957,V1125C957,V2109C957,V2205C957,C957V571,C957V728,C957V1027,C957V1125,C957V2109,C957V2205,end_cn957);
C958:CNPU6_6 port map (start_cn,clk,rst,V572C958,V729C958,V1028C958,V1126C958,V2110C958,V2206C958,C958V572,C958V729,C958V1028,C958V1126,C958V2110,C958V2206,end_cn958);
C959:CNPU6_6 port map (start_cn,clk,rst,V573C959,V730C959,V1029C959,V1127C959,V2111C959,V2207C959,C959V573,C959V730,C959V1029,C959V1127,C959V2111,C959V2207,end_cn959);
C960:CNPU6_6 port map (start_cn,clk,rst,V574C960,V731C960,V1030C960,V1128C960,V2112C960,V2208C960,C960V574,C960V731,C960V1030,C960V1128,C960V2112,C960V2208,end_cn960);
C961:CNPU6_6 port map (start_cn,clk,rst,V200C961,V354C961,V808C961,V914C961,V2113C961,V2209C961,C961V200,C961V354,C961V808,C961V914,C961V2113,C961V2209,end_cn961);
C962:CNPU6_6 port map (start_cn,clk,rst,V201C962,V355C962,V809C962,V915C962,V2114C962,V2210C962,C962V201,C962V355,C962V809,C962V915,C962V2114,C962V2210,end_cn962);
C963:CNPU6_6 port map (start_cn,clk,rst,V202C963,V356C963,V810C963,V916C963,V2115C963,V2211C963,C963V202,C963V356,C963V810,C963V916,C963V2115,C963V2211,end_cn963);
C964:CNPU6_6 port map (start_cn,clk,rst,V203C964,V357C964,V811C964,V917C964,V2116C964,V2212C964,C964V203,C964V357,C964V811,C964V917,C964V2116,C964V2212,end_cn964);
C965:CNPU6_6 port map (start_cn,clk,rst,V204C965,V358C965,V812C965,V918C965,V2117C965,V2213C965,C965V204,C965V358,C965V812,C965V918,C965V2117,C965V2213,end_cn965);
C966:CNPU6_6 port map (start_cn,clk,rst,V205C966,V359C966,V813C966,V919C966,V2118C966,V2214C966,C966V205,C966V359,C966V813,C966V919,C966V2118,C966V2214,end_cn966);
C967:CNPU6_6 port map (start_cn,clk,rst,V206C967,V360C967,V814C967,V920C967,V2119C967,V2215C967,C967V206,C967V360,C967V814,C967V920,C967V2119,C967V2215,end_cn967);
C968:CNPU6_6 port map (start_cn,clk,rst,V207C968,V361C968,V815C968,V921C968,V2120C968,V2216C968,C968V207,C968V361,C968V815,C968V921,C968V2120,C968V2216,end_cn968);
C969:CNPU6_6 port map (start_cn,clk,rst,V208C969,V362C969,V816C969,V922C969,V2121C969,V2217C969,C969V208,C969V362,C969V816,C969V922,C969V2121,C969V2217,end_cn969);
C970:CNPU6_6 port map (start_cn,clk,rst,V209C970,V363C970,V817C970,V923C970,V2122C970,V2218C970,C970V209,C970V363,C970V817,C970V923,C970V2122,C970V2218,end_cn970);
C971:CNPU6_6 port map (start_cn,clk,rst,V210C971,V364C971,V818C971,V924C971,V2123C971,V2219C971,C971V210,C971V364,C971V818,C971V924,C971V2123,C971V2219,end_cn971);
C972:CNPU6_6 port map (start_cn,clk,rst,V211C972,V365C972,V819C972,V925C972,V2124C972,V2220C972,C972V211,C972V365,C972V819,C972V925,C972V2124,C972V2220,end_cn972);
C973:CNPU6_6 port map (start_cn,clk,rst,V212C973,V366C973,V820C973,V926C973,V2125C973,V2221C973,C973V212,C973V366,C973V820,C973V926,C973V2125,C973V2221,end_cn973);
C974:CNPU6_6 port map (start_cn,clk,rst,V213C974,V367C974,V821C974,V927C974,V2126C974,V2222C974,C974V213,C974V367,C974V821,C974V927,C974V2126,C974V2222,end_cn974);
C975:CNPU6_6 port map (start_cn,clk,rst,V214C975,V368C975,V822C975,V928C975,V2127C975,V2223C975,C975V214,C975V368,C975V822,C975V928,C975V2127,C975V2223,end_cn975);
C976:CNPU6_6 port map (start_cn,clk,rst,V215C976,V369C976,V823C976,V929C976,V2128C976,V2224C976,C976V215,C976V369,C976V823,C976V929,C976V2128,C976V2224,end_cn976);
C977:CNPU6_6 port map (start_cn,clk,rst,V216C977,V370C977,V824C977,V930C977,V2129C977,V2225C977,C977V216,C977V370,C977V824,C977V930,C977V2129,C977V2225,end_cn977);
C978:CNPU6_6 port map (start_cn,clk,rst,V217C978,V371C978,V825C978,V931C978,V2130C978,V2226C978,C978V217,C978V371,C978V825,C978V931,C978V2130,C978V2226,end_cn978);
C979:CNPU6_6 port map (start_cn,clk,rst,V218C979,V372C979,V826C979,V932C979,V2131C979,V2227C979,C979V218,C979V372,C979V826,C979V932,C979V2131,C979V2227,end_cn979);
C980:CNPU6_6 port map (start_cn,clk,rst,V219C980,V373C980,V827C980,V933C980,V2132C980,V2228C980,C980V219,C980V373,C980V827,C980V933,C980V2132,C980V2228,end_cn980);
C981:CNPU6_6 port map (start_cn,clk,rst,V220C981,V374C981,V828C981,V934C981,V2133C981,V2229C981,C981V220,C981V374,C981V828,C981V934,C981V2133,C981V2229,end_cn981);
C982:CNPU6_6 port map (start_cn,clk,rst,V221C982,V375C982,V829C982,V935C982,V2134C982,V2230C982,C982V221,C982V375,C982V829,C982V935,C982V2134,C982V2230,end_cn982);
C983:CNPU6_6 port map (start_cn,clk,rst,V222C983,V376C983,V830C983,V936C983,V2135C983,V2231C983,C983V222,C983V376,C983V830,C983V936,C983V2135,C983V2231,end_cn983);
C984:CNPU6_6 port map (start_cn,clk,rst,V223C984,V377C984,V831C984,V937C984,V2136C984,V2232C984,C984V223,C984V377,C984V831,C984V937,C984V2136,C984V2232,end_cn984);
C985:CNPU6_6 port map (start_cn,clk,rst,V224C985,V378C985,V832C985,V938C985,V2137C985,V2233C985,C985V224,C985V378,C985V832,C985V938,C985V2137,C985V2233,end_cn985);
C986:CNPU6_6 port map (start_cn,clk,rst,V225C986,V379C986,V833C986,V939C986,V2138C986,V2234C986,C986V225,C986V379,C986V833,C986V939,C986V2138,C986V2234,end_cn986);
C987:CNPU6_6 port map (start_cn,clk,rst,V226C987,V380C987,V834C987,V940C987,V2139C987,V2235C987,C987V226,C987V380,C987V834,C987V940,C987V2139,C987V2235,end_cn987);
C988:CNPU6_6 port map (start_cn,clk,rst,V227C988,V381C988,V835C988,V941C988,V2140C988,V2236C988,C988V227,C988V381,C988V835,C988V941,C988V2140,C988V2236,end_cn988);
C989:CNPU6_6 port map (start_cn,clk,rst,V228C989,V382C989,V836C989,V942C989,V2141C989,V2237C989,C989V228,C989V382,C989V836,C989V942,C989V2141,C989V2237,end_cn989);
C990:CNPU6_6 port map (start_cn,clk,rst,V229C990,V383C990,V837C990,V943C990,V2142C990,V2238C990,C990V229,C990V383,C990V837,C990V943,C990V2142,C990V2238,end_cn990);
C991:CNPU6_6 port map (start_cn,clk,rst,V230C991,V384C991,V838C991,V944C991,V2143C991,V2239C991,C991V230,C991V384,C991V838,C991V944,C991V2143,C991V2239,end_cn991);
C992:CNPU6_6 port map (start_cn,clk,rst,V231C992,V289C992,V839C992,V945C992,V2144C992,V2240C992,C992V231,C992V289,C992V839,C992V945,C992V2144,C992V2240,end_cn992);
C993:CNPU6_6 port map (start_cn,clk,rst,V232C993,V290C993,V840C993,V946C993,V2145C993,V2241C993,C993V232,C993V290,C993V840,C993V946,C993V2145,C993V2241,end_cn993);
C994:CNPU6_6 port map (start_cn,clk,rst,V233C994,V291C994,V841C994,V947C994,V2146C994,V2242C994,C994V233,C994V291,C994V841,C994V947,C994V2146,C994V2242,end_cn994);
C995:CNPU6_6 port map (start_cn,clk,rst,V234C995,V292C995,V842C995,V948C995,V2147C995,V2243C995,C995V234,C995V292,C995V842,C995V948,C995V2147,C995V2243,end_cn995);
C996:CNPU6_6 port map (start_cn,clk,rst,V235C996,V293C996,V843C996,V949C996,V2148C996,V2244C996,C996V235,C996V293,C996V843,C996V949,C996V2148,C996V2244,end_cn996);
C997:CNPU6_6 port map (start_cn,clk,rst,V236C997,V294C997,V844C997,V950C997,V2149C997,V2245C997,C997V236,C997V294,C997V844,C997V950,C997V2149,C997V2245,end_cn997);
C998:CNPU6_6 port map (start_cn,clk,rst,V237C998,V295C998,V845C998,V951C998,V2150C998,V2246C998,C998V237,C998V295,C998V845,C998V951,C998V2150,C998V2246,end_cn998);
C999:CNPU6_6 port map (start_cn,clk,rst,V238C999,V296C999,V846C999,V952C999,V2151C999,V2247C999,C999V238,C999V296,C999V846,C999V952,C999V2151,C999V2247,end_cn999);
C1000:CNPU6_6 port map (start_cn,clk,rst,V239C1000,V297C1000,V847C1000,V953C1000,V2152C1000,V2248C1000,C1000V239,C1000V297,C1000V847,C1000V953,C1000V2152,C1000V2248,end_cn1000);
C1001:CNPU6_6 port map (start_cn,clk,rst,V240C1001,V298C1001,V848C1001,V954C1001,V2153C1001,V2249C1001,C1001V240,C1001V298,C1001V848,C1001V954,C1001V2153,C1001V2249,end_cn1001);
C1002:CNPU6_6 port map (start_cn,clk,rst,V241C1002,V299C1002,V849C1002,V955C1002,V2154C1002,V2250C1002,C1002V241,C1002V299,C1002V849,C1002V955,C1002V2154,C1002V2250,end_cn1002);
C1003:CNPU6_6 port map (start_cn,clk,rst,V242C1003,V300C1003,V850C1003,V956C1003,V2155C1003,V2251C1003,C1003V242,C1003V300,C1003V850,C1003V956,C1003V2155,C1003V2251,end_cn1003);
C1004:CNPU6_6 port map (start_cn,clk,rst,V243C1004,V301C1004,V851C1004,V957C1004,V2156C1004,V2252C1004,C1004V243,C1004V301,C1004V851,C1004V957,C1004V2156,C1004V2252,end_cn1004);
C1005:CNPU6_6 port map (start_cn,clk,rst,V244C1005,V302C1005,V852C1005,V958C1005,V2157C1005,V2253C1005,C1005V244,C1005V302,C1005V852,C1005V958,C1005V2157,C1005V2253,end_cn1005);
C1006:CNPU6_6 port map (start_cn,clk,rst,V245C1006,V303C1006,V853C1006,V959C1006,V2158C1006,V2254C1006,C1006V245,C1006V303,C1006V853,C1006V959,C1006V2158,C1006V2254,end_cn1006);
C1007:CNPU6_6 port map (start_cn,clk,rst,V246C1007,V304C1007,V854C1007,V960C1007,V2159C1007,V2255C1007,C1007V246,C1007V304,C1007V854,C1007V960,C1007V2159,C1007V2255,end_cn1007);
C1008:CNPU6_6 port map (start_cn,clk,rst,V247C1008,V305C1008,V855C1008,V865C1008,V2160C1008,V2256C1008,C1008V247,C1008V305,C1008V855,C1008V865,C1008V2160,C1008V2256,end_cn1008);
C1009:CNPU6_6 port map (start_cn,clk,rst,V248C1009,V306C1009,V856C1009,V866C1009,V2161C1009,V2257C1009,C1009V248,C1009V306,C1009V856,C1009V866,C1009V2161,C1009V2257,end_cn1009);
C1010:CNPU6_6 port map (start_cn,clk,rst,V249C1010,V307C1010,V857C1010,V867C1010,V2162C1010,V2258C1010,C1010V249,C1010V307,C1010V857,C1010V867,C1010V2162,C1010V2258,end_cn1010);
C1011:CNPU6_6 port map (start_cn,clk,rst,V250C1011,V308C1011,V858C1011,V868C1011,V2163C1011,V2259C1011,C1011V250,C1011V308,C1011V858,C1011V868,C1011V2163,C1011V2259,end_cn1011);
C1012:CNPU6_6 port map (start_cn,clk,rst,V251C1012,V309C1012,V859C1012,V869C1012,V2164C1012,V2260C1012,C1012V251,C1012V309,C1012V859,C1012V869,C1012V2164,C1012V2260,end_cn1012);
C1013:CNPU6_6 port map (start_cn,clk,rst,V252C1013,V310C1013,V860C1013,V870C1013,V2165C1013,V2261C1013,C1013V252,C1013V310,C1013V860,C1013V870,C1013V2165,C1013V2261,end_cn1013);
C1014:CNPU6_6 port map (start_cn,clk,rst,V253C1014,V311C1014,V861C1014,V871C1014,V2166C1014,V2262C1014,C1014V253,C1014V311,C1014V861,C1014V871,C1014V2166,C1014V2262,end_cn1014);
C1015:CNPU6_6 port map (start_cn,clk,rst,V254C1015,V312C1015,V862C1015,V872C1015,V2167C1015,V2263C1015,C1015V254,C1015V312,C1015V862,C1015V872,C1015V2167,C1015V2263,end_cn1015);
C1016:CNPU6_6 port map (start_cn,clk,rst,V255C1016,V313C1016,V863C1016,V873C1016,V2168C1016,V2264C1016,C1016V255,C1016V313,C1016V863,C1016V873,C1016V2168,C1016V2264,end_cn1016);
C1017:CNPU6_6 port map (start_cn,clk,rst,V256C1017,V314C1017,V864C1017,V874C1017,V2169C1017,V2265C1017,C1017V256,C1017V314,C1017V864,C1017V874,C1017V2169,C1017V2265,end_cn1017);
C1018:CNPU6_6 port map (start_cn,clk,rst,V257C1018,V315C1018,V769C1018,V875C1018,V2170C1018,V2266C1018,C1018V257,C1018V315,C1018V769,C1018V875,C1018V2170,C1018V2266,end_cn1018);
C1019:CNPU6_6 port map (start_cn,clk,rst,V258C1019,V316C1019,V770C1019,V876C1019,V2171C1019,V2267C1019,C1019V258,C1019V316,C1019V770,C1019V876,C1019V2171,C1019V2267,end_cn1019);
C1020:CNPU6_6 port map (start_cn,clk,rst,V259C1020,V317C1020,V771C1020,V877C1020,V2172C1020,V2268C1020,C1020V259,C1020V317,C1020V771,C1020V877,C1020V2172,C1020V2268,end_cn1020);
C1021:CNPU6_6 port map (start_cn,clk,rst,V260C1021,V318C1021,V772C1021,V878C1021,V2173C1021,V2269C1021,C1021V260,C1021V318,C1021V772,C1021V878,C1021V2173,C1021V2269,end_cn1021);
C1022:CNPU6_6 port map (start_cn,clk,rst,V261C1022,V319C1022,V773C1022,V879C1022,V2174C1022,V2270C1022,C1022V261,C1022V319,C1022V773,C1022V879,C1022V2174,C1022V2270,end_cn1022);
C1023:CNPU6_6 port map (start_cn,clk,rst,V262C1023,V320C1023,V774C1023,V880C1023,V2175C1023,V2271C1023,C1023V262,C1023V320,C1023V774,C1023V880,C1023V2175,C1023V2271,end_cn1023);
C1024:CNPU6_6 port map (start_cn,clk,rst,V263C1024,V321C1024,V775C1024,V881C1024,V2176C1024,V2272C1024,C1024V263,C1024V321,C1024V775,C1024V881,C1024V2176,C1024V2272,end_cn1024);
C1025:CNPU6_6 port map (start_cn,clk,rst,V264C1025,V322C1025,V776C1025,V882C1025,V2177C1025,V2273C1025,C1025V264,C1025V322,C1025V776,C1025V882,C1025V2177,C1025V2273,end_cn1025);
C1026:CNPU6_6 port map (start_cn,clk,rst,V265C1026,V323C1026,V777C1026,V883C1026,V2178C1026,V2274C1026,C1026V265,C1026V323,C1026V777,C1026V883,C1026V2178,C1026V2274,end_cn1026);
C1027:CNPU6_6 port map (start_cn,clk,rst,V266C1027,V324C1027,V778C1027,V884C1027,V2179C1027,V2275C1027,C1027V266,C1027V324,C1027V778,C1027V884,C1027V2179,C1027V2275,end_cn1027);
C1028:CNPU6_6 port map (start_cn,clk,rst,V267C1028,V325C1028,V779C1028,V885C1028,V2180C1028,V2276C1028,C1028V267,C1028V325,C1028V779,C1028V885,C1028V2180,C1028V2276,end_cn1028);
C1029:CNPU6_6 port map (start_cn,clk,rst,V268C1029,V326C1029,V780C1029,V886C1029,V2181C1029,V2277C1029,C1029V268,C1029V326,C1029V780,C1029V886,C1029V2181,C1029V2277,end_cn1029);
C1030:CNPU6_6 port map (start_cn,clk,rst,V269C1030,V327C1030,V781C1030,V887C1030,V2182C1030,V2278C1030,C1030V269,C1030V327,C1030V781,C1030V887,C1030V2182,C1030V2278,end_cn1030);
C1031:CNPU6_6 port map (start_cn,clk,rst,V270C1031,V328C1031,V782C1031,V888C1031,V2183C1031,V2279C1031,C1031V270,C1031V328,C1031V782,C1031V888,C1031V2183,C1031V2279,end_cn1031);
C1032:CNPU6_6 port map (start_cn,clk,rst,V271C1032,V329C1032,V783C1032,V889C1032,V2184C1032,V2280C1032,C1032V271,C1032V329,C1032V783,C1032V889,C1032V2184,C1032V2280,end_cn1032);
C1033:CNPU6_6 port map (start_cn,clk,rst,V272C1033,V330C1033,V784C1033,V890C1033,V2185C1033,V2281C1033,C1033V272,C1033V330,C1033V784,C1033V890,C1033V2185,C1033V2281,end_cn1033);
C1034:CNPU6_6 port map (start_cn,clk,rst,V273C1034,V331C1034,V785C1034,V891C1034,V2186C1034,V2282C1034,C1034V273,C1034V331,C1034V785,C1034V891,C1034V2186,C1034V2282,end_cn1034);
C1035:CNPU6_6 port map (start_cn,clk,rst,V274C1035,V332C1035,V786C1035,V892C1035,V2187C1035,V2283C1035,C1035V274,C1035V332,C1035V786,C1035V892,C1035V2187,C1035V2283,end_cn1035);
C1036:CNPU6_6 port map (start_cn,clk,rst,V275C1036,V333C1036,V787C1036,V893C1036,V2188C1036,V2284C1036,C1036V275,C1036V333,C1036V787,C1036V893,C1036V2188,C1036V2284,end_cn1036);
C1037:CNPU6_6 port map (start_cn,clk,rst,V276C1037,V334C1037,V788C1037,V894C1037,V2189C1037,V2285C1037,C1037V276,C1037V334,C1037V788,C1037V894,C1037V2189,C1037V2285,end_cn1037);
C1038:CNPU6_6 port map (start_cn,clk,rst,V277C1038,V335C1038,V789C1038,V895C1038,V2190C1038,V2286C1038,C1038V277,C1038V335,C1038V789,C1038V895,C1038V2190,C1038V2286,end_cn1038);
C1039:CNPU6_6 port map (start_cn,clk,rst,V278C1039,V336C1039,V790C1039,V896C1039,V2191C1039,V2287C1039,C1039V278,C1039V336,C1039V790,C1039V896,C1039V2191,C1039V2287,end_cn1039);
C1040:CNPU6_6 port map (start_cn,clk,rst,V279C1040,V337C1040,V791C1040,V897C1040,V2192C1040,V2288C1040,C1040V279,C1040V337,C1040V791,C1040V897,C1040V2192,C1040V2288,end_cn1040);
C1041:CNPU6_6 port map (start_cn,clk,rst,V280C1041,V338C1041,V792C1041,V898C1041,V2193C1041,V2289C1041,C1041V280,C1041V338,C1041V792,C1041V898,C1041V2193,C1041V2289,end_cn1041);
C1042:CNPU6_6 port map (start_cn,clk,rst,V281C1042,V339C1042,V793C1042,V899C1042,V2194C1042,V2290C1042,C1042V281,C1042V339,C1042V793,C1042V899,C1042V2194,C1042V2290,end_cn1042);
C1043:CNPU6_6 port map (start_cn,clk,rst,V282C1043,V340C1043,V794C1043,V900C1043,V2195C1043,V2291C1043,C1043V282,C1043V340,C1043V794,C1043V900,C1043V2195,C1043V2291,end_cn1043);
C1044:CNPU6_6 port map (start_cn,clk,rst,V283C1044,V341C1044,V795C1044,V901C1044,V2196C1044,V2292C1044,C1044V283,C1044V341,C1044V795,C1044V901,C1044V2196,C1044V2292,end_cn1044);
C1045:CNPU6_6 port map (start_cn,clk,rst,V284C1045,V342C1045,V796C1045,V902C1045,V2197C1045,V2293C1045,C1045V284,C1045V342,C1045V796,C1045V902,C1045V2197,C1045V2293,end_cn1045);
C1046:CNPU6_6 port map (start_cn,clk,rst,V285C1046,V343C1046,V797C1046,V903C1046,V2198C1046,V2294C1046,C1046V285,C1046V343,C1046V797,C1046V903,C1046V2198,C1046V2294,end_cn1046);
C1047:CNPU6_6 port map (start_cn,clk,rst,V286C1047,V344C1047,V798C1047,V904C1047,V2199C1047,V2295C1047,C1047V286,C1047V344,C1047V798,C1047V904,C1047V2199,C1047V2295,end_cn1047);
C1048:CNPU6_6 port map (start_cn,clk,rst,V287C1048,V345C1048,V799C1048,V905C1048,V2200C1048,V2296C1048,C1048V287,C1048V345,C1048V799,C1048V905,C1048V2200,C1048V2296,end_cn1048);
C1049:CNPU6_6 port map (start_cn,clk,rst,V288C1049,V346C1049,V800C1049,V906C1049,V2201C1049,V2297C1049,C1049V288,C1049V346,C1049V800,C1049V906,C1049V2201,C1049V2297,end_cn1049);
C1050:CNPU6_6 port map (start_cn,clk,rst,V193C1050,V347C1050,V801C1050,V907C1050,V2202C1050,V2298C1050,C1050V193,C1050V347,C1050V801,C1050V907,C1050V2202,C1050V2298,end_cn1050);
C1051:CNPU6_6 port map (start_cn,clk,rst,V194C1051,V348C1051,V802C1051,V908C1051,V2203C1051,V2299C1051,C1051V194,C1051V348,C1051V802,C1051V908,C1051V2203,C1051V2299,end_cn1051);
C1052:CNPU6_6 port map (start_cn,clk,rst,V195C1052,V349C1052,V803C1052,V909C1052,V2204C1052,V2300C1052,C1052V195,C1052V349,C1052V803,C1052V909,C1052V2204,C1052V2300,end_cn1052);
C1053:CNPU6_6 port map (start_cn,clk,rst,V196C1053,V350C1053,V804C1053,V910C1053,V2205C1053,V2301C1053,C1053V196,C1053V350,C1053V804,C1053V910,C1053V2205,C1053V2301,end_cn1053);
C1054:CNPU6_6 port map (start_cn,clk,rst,V197C1054,V351C1054,V805C1054,V911C1054,V2206C1054,V2302C1054,C1054V197,C1054V351,C1054V805,C1054V911,C1054V2206,C1054V2302,end_cn1054);
C1055:CNPU6_6 port map (start_cn,clk,rst,V198C1055,V352C1055,V806C1055,V912C1055,V2207C1055,V2303C1055,C1055V198,C1055V352,C1055V806,C1055V912,C1055V2207,C1055V2303,end_cn1055);
C1056:CNPU6_6 port map (start_cn,clk,rst,V199C1056,V353C1056,V807C1056,V913C1056,V2208C1056,V2304C1056,C1056V199,C1056V353,C1056V807,C1056V913,C1056V2208,C1056V2304,end_cn1056);
C1057:CNPU6_6 port map (start_cn,clk,rst,V44C1057,V547C1057,V714C1057,V1083C1057,V1160C1057,V2209C1057,C1057V44,C1057V547,C1057V714,C1057V1083,C1057V1160,C1057V2209,end_cn1057);
C1058:CNPU6_6 port map (start_cn,clk,rst,V45C1058,V548C1058,V715C1058,V1084C1058,V1161C1058,V2210C1058,C1058V45,C1058V548,C1058V715,C1058V1084,C1058V1161,C1058V2210,end_cn1058);
C1059:CNPU6_6 port map (start_cn,clk,rst,V46C1059,V549C1059,V716C1059,V1085C1059,V1162C1059,V2211C1059,C1059V46,C1059V549,C1059V716,C1059V1085,C1059V1162,C1059V2211,end_cn1059);
C1060:CNPU6_6 port map (start_cn,clk,rst,V47C1060,V550C1060,V717C1060,V1086C1060,V1163C1060,V2212C1060,C1060V47,C1060V550,C1060V717,C1060V1086,C1060V1163,C1060V2212,end_cn1060);
C1061:CNPU6_6 port map (start_cn,clk,rst,V48C1061,V551C1061,V718C1061,V1087C1061,V1164C1061,V2213C1061,C1061V48,C1061V551,C1061V718,C1061V1087,C1061V1164,C1061V2213,end_cn1061);
C1062:CNPU6_6 port map (start_cn,clk,rst,V49C1062,V552C1062,V719C1062,V1088C1062,V1165C1062,V2214C1062,C1062V49,C1062V552,C1062V719,C1062V1088,C1062V1165,C1062V2214,end_cn1062);
C1063:CNPU6_6 port map (start_cn,clk,rst,V50C1063,V553C1063,V720C1063,V1089C1063,V1166C1063,V2215C1063,C1063V50,C1063V553,C1063V720,C1063V1089,C1063V1166,C1063V2215,end_cn1063);
C1064:CNPU6_6 port map (start_cn,clk,rst,V51C1064,V554C1064,V721C1064,V1090C1064,V1167C1064,V2216C1064,C1064V51,C1064V554,C1064V721,C1064V1090,C1064V1167,C1064V2216,end_cn1064);
C1065:CNPU6_6 port map (start_cn,clk,rst,V52C1065,V555C1065,V722C1065,V1091C1065,V1168C1065,V2217C1065,C1065V52,C1065V555,C1065V722,C1065V1091,C1065V1168,C1065V2217,end_cn1065);
C1066:CNPU6_6 port map (start_cn,clk,rst,V53C1066,V556C1066,V723C1066,V1092C1066,V1169C1066,V2218C1066,C1066V53,C1066V556,C1066V723,C1066V1092,C1066V1169,C1066V2218,end_cn1066);
C1067:CNPU6_6 port map (start_cn,clk,rst,V54C1067,V557C1067,V724C1067,V1093C1067,V1170C1067,V2219C1067,C1067V54,C1067V557,C1067V724,C1067V1093,C1067V1170,C1067V2219,end_cn1067);
C1068:CNPU6_6 port map (start_cn,clk,rst,V55C1068,V558C1068,V725C1068,V1094C1068,V1171C1068,V2220C1068,C1068V55,C1068V558,C1068V725,C1068V1094,C1068V1171,C1068V2220,end_cn1068);
C1069:CNPU6_6 port map (start_cn,clk,rst,V56C1069,V559C1069,V726C1069,V1095C1069,V1172C1069,V2221C1069,C1069V56,C1069V559,C1069V726,C1069V1095,C1069V1172,C1069V2221,end_cn1069);
C1070:CNPU6_6 port map (start_cn,clk,rst,V57C1070,V560C1070,V727C1070,V1096C1070,V1173C1070,V2222C1070,C1070V57,C1070V560,C1070V727,C1070V1096,C1070V1173,C1070V2222,end_cn1070);
C1071:CNPU6_6 port map (start_cn,clk,rst,V58C1071,V561C1071,V728C1071,V1097C1071,V1174C1071,V2223C1071,C1071V58,C1071V561,C1071V728,C1071V1097,C1071V1174,C1071V2223,end_cn1071);
C1072:CNPU6_6 port map (start_cn,clk,rst,V59C1072,V562C1072,V729C1072,V1098C1072,V1175C1072,V2224C1072,C1072V59,C1072V562,C1072V729,C1072V1098,C1072V1175,C1072V2224,end_cn1072);
C1073:CNPU6_6 port map (start_cn,clk,rst,V60C1073,V563C1073,V730C1073,V1099C1073,V1176C1073,V2225C1073,C1073V60,C1073V563,C1073V730,C1073V1099,C1073V1176,C1073V2225,end_cn1073);
C1074:CNPU6_6 port map (start_cn,clk,rst,V61C1074,V564C1074,V731C1074,V1100C1074,V1177C1074,V2226C1074,C1074V61,C1074V564,C1074V731,C1074V1100,C1074V1177,C1074V2226,end_cn1074);
C1075:CNPU6_6 port map (start_cn,clk,rst,V62C1075,V565C1075,V732C1075,V1101C1075,V1178C1075,V2227C1075,C1075V62,C1075V565,C1075V732,C1075V1101,C1075V1178,C1075V2227,end_cn1075);
C1076:CNPU6_6 port map (start_cn,clk,rst,V63C1076,V566C1076,V733C1076,V1102C1076,V1179C1076,V2228C1076,C1076V63,C1076V566,C1076V733,C1076V1102,C1076V1179,C1076V2228,end_cn1076);
C1077:CNPU6_6 port map (start_cn,clk,rst,V64C1077,V567C1077,V734C1077,V1103C1077,V1180C1077,V2229C1077,C1077V64,C1077V567,C1077V734,C1077V1103,C1077V1180,C1077V2229,end_cn1077);
C1078:CNPU6_6 port map (start_cn,clk,rst,V65C1078,V568C1078,V735C1078,V1104C1078,V1181C1078,V2230C1078,C1078V65,C1078V568,C1078V735,C1078V1104,C1078V1181,C1078V2230,end_cn1078);
C1079:CNPU6_6 port map (start_cn,clk,rst,V66C1079,V569C1079,V736C1079,V1105C1079,V1182C1079,V2231C1079,C1079V66,C1079V569,C1079V736,C1079V1105,C1079V1182,C1079V2231,end_cn1079);
C1080:CNPU6_6 port map (start_cn,clk,rst,V67C1080,V570C1080,V737C1080,V1106C1080,V1183C1080,V2232C1080,C1080V67,C1080V570,C1080V737,C1080V1106,C1080V1183,C1080V2232,end_cn1080);
C1081:CNPU6_6 port map (start_cn,clk,rst,V68C1081,V571C1081,V738C1081,V1107C1081,V1184C1081,V2233C1081,C1081V68,C1081V571,C1081V738,C1081V1107,C1081V1184,C1081V2233,end_cn1081);
C1082:CNPU6_6 port map (start_cn,clk,rst,V69C1082,V572C1082,V739C1082,V1108C1082,V1185C1082,V2234C1082,C1082V69,C1082V572,C1082V739,C1082V1108,C1082V1185,C1082V2234,end_cn1082);
C1083:CNPU6_6 port map (start_cn,clk,rst,V70C1083,V573C1083,V740C1083,V1109C1083,V1186C1083,V2235C1083,C1083V70,C1083V573,C1083V740,C1083V1109,C1083V1186,C1083V2235,end_cn1083);
C1084:CNPU6_6 port map (start_cn,clk,rst,V71C1084,V574C1084,V741C1084,V1110C1084,V1187C1084,V2236C1084,C1084V71,C1084V574,C1084V741,C1084V1110,C1084V1187,C1084V2236,end_cn1084);
C1085:CNPU6_6 port map (start_cn,clk,rst,V72C1085,V575C1085,V742C1085,V1111C1085,V1188C1085,V2237C1085,C1085V72,C1085V575,C1085V742,C1085V1111,C1085V1188,C1085V2237,end_cn1085);
C1086:CNPU6_6 port map (start_cn,clk,rst,V73C1086,V576C1086,V743C1086,V1112C1086,V1189C1086,V2238C1086,C1086V73,C1086V576,C1086V743,C1086V1112,C1086V1189,C1086V2238,end_cn1086);
C1087:CNPU6_6 port map (start_cn,clk,rst,V74C1087,V481C1087,V744C1087,V1113C1087,V1190C1087,V2239C1087,C1087V74,C1087V481,C1087V744,C1087V1113,C1087V1190,C1087V2239,end_cn1087);
C1088:CNPU6_6 port map (start_cn,clk,rst,V75C1088,V482C1088,V745C1088,V1114C1088,V1191C1088,V2240C1088,C1088V75,C1088V482,C1088V745,C1088V1114,C1088V1191,C1088V2240,end_cn1088);
C1089:CNPU6_6 port map (start_cn,clk,rst,V76C1089,V483C1089,V746C1089,V1115C1089,V1192C1089,V2241C1089,C1089V76,C1089V483,C1089V746,C1089V1115,C1089V1192,C1089V2241,end_cn1089);
C1090:CNPU6_6 port map (start_cn,clk,rst,V77C1090,V484C1090,V747C1090,V1116C1090,V1193C1090,V2242C1090,C1090V77,C1090V484,C1090V747,C1090V1116,C1090V1193,C1090V2242,end_cn1090);
C1091:CNPU6_6 port map (start_cn,clk,rst,V78C1091,V485C1091,V748C1091,V1117C1091,V1194C1091,V2243C1091,C1091V78,C1091V485,C1091V748,C1091V1117,C1091V1194,C1091V2243,end_cn1091);
C1092:CNPU6_6 port map (start_cn,clk,rst,V79C1092,V486C1092,V749C1092,V1118C1092,V1195C1092,V2244C1092,C1092V79,C1092V486,C1092V749,C1092V1118,C1092V1195,C1092V2244,end_cn1092);
C1093:CNPU6_6 port map (start_cn,clk,rst,V80C1093,V487C1093,V750C1093,V1119C1093,V1196C1093,V2245C1093,C1093V80,C1093V487,C1093V750,C1093V1119,C1093V1196,C1093V2245,end_cn1093);
C1094:CNPU6_6 port map (start_cn,clk,rst,V81C1094,V488C1094,V751C1094,V1120C1094,V1197C1094,V2246C1094,C1094V81,C1094V488,C1094V751,C1094V1120,C1094V1197,C1094V2246,end_cn1094);
C1095:CNPU6_6 port map (start_cn,clk,rst,V82C1095,V489C1095,V752C1095,V1121C1095,V1198C1095,V2247C1095,C1095V82,C1095V489,C1095V752,C1095V1121,C1095V1198,C1095V2247,end_cn1095);
C1096:CNPU6_6 port map (start_cn,clk,rst,V83C1096,V490C1096,V753C1096,V1122C1096,V1199C1096,V2248C1096,C1096V83,C1096V490,C1096V753,C1096V1122,C1096V1199,C1096V2248,end_cn1096);
C1097:CNPU6_6 port map (start_cn,clk,rst,V84C1097,V491C1097,V754C1097,V1123C1097,V1200C1097,V2249C1097,C1097V84,C1097V491,C1097V754,C1097V1123,C1097V1200,C1097V2249,end_cn1097);
C1098:CNPU6_6 port map (start_cn,clk,rst,V85C1098,V492C1098,V755C1098,V1124C1098,V1201C1098,V2250C1098,C1098V85,C1098V492,C1098V755,C1098V1124,C1098V1201,C1098V2250,end_cn1098);
C1099:CNPU6_6 port map (start_cn,clk,rst,V86C1099,V493C1099,V756C1099,V1125C1099,V1202C1099,V2251C1099,C1099V86,C1099V493,C1099V756,C1099V1125,C1099V1202,C1099V2251,end_cn1099);
C1100:CNPU6_6 port map (start_cn,clk,rst,V87C1100,V494C1100,V757C1100,V1126C1100,V1203C1100,V2252C1100,C1100V87,C1100V494,C1100V757,C1100V1126,C1100V1203,C1100V2252,end_cn1100);
C1101:CNPU6_6 port map (start_cn,clk,rst,V88C1101,V495C1101,V758C1101,V1127C1101,V1204C1101,V2253C1101,C1101V88,C1101V495,C1101V758,C1101V1127,C1101V1204,C1101V2253,end_cn1101);
C1102:CNPU6_6 port map (start_cn,clk,rst,V89C1102,V496C1102,V759C1102,V1128C1102,V1205C1102,V2254C1102,C1102V89,C1102V496,C1102V759,C1102V1128,C1102V1205,C1102V2254,end_cn1102);
C1103:CNPU6_6 port map (start_cn,clk,rst,V90C1103,V497C1103,V760C1103,V1129C1103,V1206C1103,V2255C1103,C1103V90,C1103V497,C1103V760,C1103V1129,C1103V1206,C1103V2255,end_cn1103);
C1104:CNPU6_6 port map (start_cn,clk,rst,V91C1104,V498C1104,V761C1104,V1130C1104,V1207C1104,V2256C1104,C1104V91,C1104V498,C1104V761,C1104V1130,C1104V1207,C1104V2256,end_cn1104);
C1105:CNPU6_6 port map (start_cn,clk,rst,V92C1105,V499C1105,V762C1105,V1131C1105,V1208C1105,V2257C1105,C1105V92,C1105V499,C1105V762,C1105V1131,C1105V1208,C1105V2257,end_cn1105);
C1106:CNPU6_6 port map (start_cn,clk,rst,V93C1106,V500C1106,V763C1106,V1132C1106,V1209C1106,V2258C1106,C1106V93,C1106V500,C1106V763,C1106V1132,C1106V1209,C1106V2258,end_cn1106);
C1107:CNPU6_6 port map (start_cn,clk,rst,V94C1107,V501C1107,V764C1107,V1133C1107,V1210C1107,V2259C1107,C1107V94,C1107V501,C1107V764,C1107V1133,C1107V1210,C1107V2259,end_cn1107);
C1108:CNPU6_6 port map (start_cn,clk,rst,V95C1108,V502C1108,V765C1108,V1134C1108,V1211C1108,V2260C1108,C1108V95,C1108V502,C1108V765,C1108V1134,C1108V1211,C1108V2260,end_cn1108);
C1109:CNPU6_6 port map (start_cn,clk,rst,V96C1109,V503C1109,V766C1109,V1135C1109,V1212C1109,V2261C1109,C1109V96,C1109V503,C1109V766,C1109V1135,C1109V1212,C1109V2261,end_cn1109);
C1110:CNPU6_6 port map (start_cn,clk,rst,V1C1110,V504C1110,V767C1110,V1136C1110,V1213C1110,V2262C1110,C1110V1,C1110V504,C1110V767,C1110V1136,C1110V1213,C1110V2262,end_cn1110);
C1111:CNPU6_6 port map (start_cn,clk,rst,V2C1111,V505C1111,V768C1111,V1137C1111,V1214C1111,V2263C1111,C1111V2,C1111V505,C1111V768,C1111V1137,C1111V1214,C1111V2263,end_cn1111);
C1112:CNPU6_6 port map (start_cn,clk,rst,V3C1112,V506C1112,V673C1112,V1138C1112,V1215C1112,V2264C1112,C1112V3,C1112V506,C1112V673,C1112V1138,C1112V1215,C1112V2264,end_cn1112);
C1113:CNPU6_6 port map (start_cn,clk,rst,V4C1113,V507C1113,V674C1113,V1139C1113,V1216C1113,V2265C1113,C1113V4,C1113V507,C1113V674,C1113V1139,C1113V1216,C1113V2265,end_cn1113);
C1114:CNPU6_6 port map (start_cn,clk,rst,V5C1114,V508C1114,V675C1114,V1140C1114,V1217C1114,V2266C1114,C1114V5,C1114V508,C1114V675,C1114V1140,C1114V1217,C1114V2266,end_cn1114);
C1115:CNPU6_6 port map (start_cn,clk,rst,V6C1115,V509C1115,V676C1115,V1141C1115,V1218C1115,V2267C1115,C1115V6,C1115V509,C1115V676,C1115V1141,C1115V1218,C1115V2267,end_cn1115);
C1116:CNPU6_6 port map (start_cn,clk,rst,V7C1116,V510C1116,V677C1116,V1142C1116,V1219C1116,V2268C1116,C1116V7,C1116V510,C1116V677,C1116V1142,C1116V1219,C1116V2268,end_cn1116);
C1117:CNPU6_6 port map (start_cn,clk,rst,V8C1117,V511C1117,V678C1117,V1143C1117,V1220C1117,V2269C1117,C1117V8,C1117V511,C1117V678,C1117V1143,C1117V1220,C1117V2269,end_cn1117);
C1118:CNPU6_6 port map (start_cn,clk,rst,V9C1118,V512C1118,V679C1118,V1144C1118,V1221C1118,V2270C1118,C1118V9,C1118V512,C1118V679,C1118V1144,C1118V1221,C1118V2270,end_cn1118);
C1119:CNPU6_6 port map (start_cn,clk,rst,V10C1119,V513C1119,V680C1119,V1145C1119,V1222C1119,V2271C1119,C1119V10,C1119V513,C1119V680,C1119V1145,C1119V1222,C1119V2271,end_cn1119);
C1120:CNPU6_6 port map (start_cn,clk,rst,V11C1120,V514C1120,V681C1120,V1146C1120,V1223C1120,V2272C1120,C1120V11,C1120V514,C1120V681,C1120V1146,C1120V1223,C1120V2272,end_cn1120);
C1121:CNPU6_6 port map (start_cn,clk,rst,V12C1121,V515C1121,V682C1121,V1147C1121,V1224C1121,V2273C1121,C1121V12,C1121V515,C1121V682,C1121V1147,C1121V1224,C1121V2273,end_cn1121);
C1122:CNPU6_6 port map (start_cn,clk,rst,V13C1122,V516C1122,V683C1122,V1148C1122,V1225C1122,V2274C1122,C1122V13,C1122V516,C1122V683,C1122V1148,C1122V1225,C1122V2274,end_cn1122);
C1123:CNPU6_6 port map (start_cn,clk,rst,V14C1123,V517C1123,V684C1123,V1149C1123,V1226C1123,V2275C1123,C1123V14,C1123V517,C1123V684,C1123V1149,C1123V1226,C1123V2275,end_cn1123);
C1124:CNPU6_6 port map (start_cn,clk,rst,V15C1124,V518C1124,V685C1124,V1150C1124,V1227C1124,V2276C1124,C1124V15,C1124V518,C1124V685,C1124V1150,C1124V1227,C1124V2276,end_cn1124);
C1125:CNPU6_6 port map (start_cn,clk,rst,V16C1125,V519C1125,V686C1125,V1151C1125,V1228C1125,V2277C1125,C1125V16,C1125V519,C1125V686,C1125V1151,C1125V1228,C1125V2277,end_cn1125);
C1126:CNPU6_6 port map (start_cn,clk,rst,V17C1126,V520C1126,V687C1126,V1152C1126,V1229C1126,V2278C1126,C1126V17,C1126V520,C1126V687,C1126V1152,C1126V1229,C1126V2278,end_cn1126);
C1127:CNPU6_6 port map (start_cn,clk,rst,V18C1127,V521C1127,V688C1127,V1057C1127,V1230C1127,V2279C1127,C1127V18,C1127V521,C1127V688,C1127V1057,C1127V1230,C1127V2279,end_cn1127);
C1128:CNPU6_6 port map (start_cn,clk,rst,V19C1128,V522C1128,V689C1128,V1058C1128,V1231C1128,V2280C1128,C1128V19,C1128V522,C1128V689,C1128V1058,C1128V1231,C1128V2280,end_cn1128);
C1129:CNPU6_6 port map (start_cn,clk,rst,V20C1129,V523C1129,V690C1129,V1059C1129,V1232C1129,V2281C1129,C1129V20,C1129V523,C1129V690,C1129V1059,C1129V1232,C1129V2281,end_cn1129);
C1130:CNPU6_6 port map (start_cn,clk,rst,V21C1130,V524C1130,V691C1130,V1060C1130,V1233C1130,V2282C1130,C1130V21,C1130V524,C1130V691,C1130V1060,C1130V1233,C1130V2282,end_cn1130);
C1131:CNPU6_6 port map (start_cn,clk,rst,V22C1131,V525C1131,V692C1131,V1061C1131,V1234C1131,V2283C1131,C1131V22,C1131V525,C1131V692,C1131V1061,C1131V1234,C1131V2283,end_cn1131);
C1132:CNPU6_6 port map (start_cn,clk,rst,V23C1132,V526C1132,V693C1132,V1062C1132,V1235C1132,V2284C1132,C1132V23,C1132V526,C1132V693,C1132V1062,C1132V1235,C1132V2284,end_cn1132);
C1133:CNPU6_6 port map (start_cn,clk,rst,V24C1133,V527C1133,V694C1133,V1063C1133,V1236C1133,V2285C1133,C1133V24,C1133V527,C1133V694,C1133V1063,C1133V1236,C1133V2285,end_cn1133);
C1134:CNPU6_6 port map (start_cn,clk,rst,V25C1134,V528C1134,V695C1134,V1064C1134,V1237C1134,V2286C1134,C1134V25,C1134V528,C1134V695,C1134V1064,C1134V1237,C1134V2286,end_cn1134);
C1135:CNPU6_6 port map (start_cn,clk,rst,V26C1135,V529C1135,V696C1135,V1065C1135,V1238C1135,V2287C1135,C1135V26,C1135V529,C1135V696,C1135V1065,C1135V1238,C1135V2287,end_cn1135);
C1136:CNPU6_6 port map (start_cn,clk,rst,V27C1136,V530C1136,V697C1136,V1066C1136,V1239C1136,V2288C1136,C1136V27,C1136V530,C1136V697,C1136V1066,C1136V1239,C1136V2288,end_cn1136);
C1137:CNPU6_6 port map (start_cn,clk,rst,V28C1137,V531C1137,V698C1137,V1067C1137,V1240C1137,V2289C1137,C1137V28,C1137V531,C1137V698,C1137V1067,C1137V1240,C1137V2289,end_cn1137);
C1138:CNPU6_6 port map (start_cn,clk,rst,V29C1138,V532C1138,V699C1138,V1068C1138,V1241C1138,V2290C1138,C1138V29,C1138V532,C1138V699,C1138V1068,C1138V1241,C1138V2290,end_cn1138);
C1139:CNPU6_6 port map (start_cn,clk,rst,V30C1139,V533C1139,V700C1139,V1069C1139,V1242C1139,V2291C1139,C1139V30,C1139V533,C1139V700,C1139V1069,C1139V1242,C1139V2291,end_cn1139);
C1140:CNPU6_6 port map (start_cn,clk,rst,V31C1140,V534C1140,V701C1140,V1070C1140,V1243C1140,V2292C1140,C1140V31,C1140V534,C1140V701,C1140V1070,C1140V1243,C1140V2292,end_cn1140);
C1141:CNPU6_6 port map (start_cn,clk,rst,V32C1141,V535C1141,V702C1141,V1071C1141,V1244C1141,V2293C1141,C1141V32,C1141V535,C1141V702,C1141V1071,C1141V1244,C1141V2293,end_cn1141);
C1142:CNPU6_6 port map (start_cn,clk,rst,V33C1142,V536C1142,V703C1142,V1072C1142,V1245C1142,V2294C1142,C1142V33,C1142V536,C1142V703,C1142V1072,C1142V1245,C1142V2294,end_cn1142);
C1143:CNPU6_6 port map (start_cn,clk,rst,V34C1143,V537C1143,V704C1143,V1073C1143,V1246C1143,V2295C1143,C1143V34,C1143V537,C1143V704,C1143V1073,C1143V1246,C1143V2295,end_cn1143);
C1144:CNPU6_6 port map (start_cn,clk,rst,V35C1144,V538C1144,V705C1144,V1074C1144,V1247C1144,V2296C1144,C1144V35,C1144V538,C1144V705,C1144V1074,C1144V1247,C1144V2296,end_cn1144);
C1145:CNPU6_6 port map (start_cn,clk,rst,V36C1145,V539C1145,V706C1145,V1075C1145,V1248C1145,V2297C1145,C1145V36,C1145V539,C1145V706,C1145V1075,C1145V1248,C1145V2297,end_cn1145);
C1146:CNPU6_6 port map (start_cn,clk,rst,V37C1146,V540C1146,V707C1146,V1076C1146,V1153C1146,V2298C1146,C1146V37,C1146V540,C1146V707,C1146V1076,C1146V1153,C1146V2298,end_cn1146);
C1147:CNPU6_6 port map (start_cn,clk,rst,V38C1147,V541C1147,V708C1147,V1077C1147,V1154C1147,V2299C1147,C1147V38,C1147V541,C1147V708,C1147V1077,C1147V1154,C1147V2299,end_cn1147);
C1148:CNPU6_6 port map (start_cn,clk,rst,V39C1148,V542C1148,V709C1148,V1078C1148,V1155C1148,V2300C1148,C1148V39,C1148V542,C1148V709,C1148V1078,C1148V1155,C1148V2300,end_cn1148);
C1149:CNPU6_6 port map (start_cn,clk,rst,V40C1149,V543C1149,V710C1149,V1079C1149,V1156C1149,V2301C1149,C1149V40,C1149V543,C1149V710,C1149V1079,C1149V1156,C1149V2301,end_cn1149);
C1150:CNPU6_6 port map (start_cn,clk,rst,V41C1150,V544C1150,V711C1150,V1080C1150,V1157C1150,V2302C1150,C1150V41,C1150V544,C1150V711,C1150V1080,C1150V1157,C1150V2302,end_cn1150);
C1151:CNPU6_6 port map (start_cn,clk,rst,V42C1151,V545C1151,V712C1151,V1081C1151,V1158C1151,V2303C1151,C1151V42,C1151V545,C1151V712,C1151V1081,C1151V1158,C1151V2303,end_cn1151);
C1152:CNPU6_6 port map (start_cn,clk,rst,V43C1152,V546C1152,V713C1152,V1082C1152,V1159C1152,V2304C1152,C1152V43,C1152V546,C1152V713,C1152V1082,C1152V1159,C1152V2304,end_cn1152);

V1:VNPU3_3 port map (start_vn,clk,rst,Lc1,C324V1,C853V1,C1110V1,V1C324,V1C853,V1C1110,SI1,end_vn1);
V2:VNPU3_3 port map (start_vn,clk,rst,Lc2,C325V2,C854V2,C1111V2,V2C325,V2C854,V2C1111,SI2,end_vn2);
V3:VNPU3_3 port map (start_vn,clk,rst,Lc3,C326V3,C855V3,C1112V3,V3C326,V3C855,V3C1112,SI3,end_vn3);
V4:VNPU3_3 port map (start_vn,clk,rst,Lc4,C327V4,C856V4,C1113V4,V4C327,V4C856,V4C1113,SI4,end_vn4);
V5:VNPU3_3 port map (start_vn,clk,rst,Lc5,C328V5,C857V5,C1114V5,V5C328,V5C857,V5C1114,SI5,end_vn5);
V6:VNPU3_3 port map (start_vn,clk,rst,Lc6,C329V6,C858V6,C1115V6,V6C329,V6C858,V6C1115,SI6,end_vn6);
V7:VNPU3_3 port map (start_vn,clk,rst,Lc7,C330V7,C859V7,C1116V7,V7C330,V7C859,V7C1116,SI7,end_vn7);
V8:VNPU3_3 port map (start_vn,clk,rst,Lc8,C331V8,C860V8,C1117V8,V8C331,V8C860,V8C1117,SI8,end_vn8);
V9:VNPU3_3 port map (start_vn,clk,rst,Lc9,C332V9,C861V9,C1118V9,V9C332,V9C861,V9C1118,SI9,end_vn9);
V10:VNPU3_3 port map (start_vn,clk,rst,Lc10,C333V10,C862V10,C1119V10,V10C333,V10C862,V10C1119,SI10,end_vn10);
V11:VNPU3_3 port map (start_vn,clk,rst,Lc11,C334V11,C863V11,C1120V11,V11C334,V11C863,V11C1120,SI11,end_vn11);
V12:VNPU3_3 port map (start_vn,clk,rst,Lc12,C335V12,C864V12,C1121V12,V12C335,V12C864,V12C1121,SI12,end_vn12);
V13:VNPU3_3 port map (start_vn,clk,rst,Lc13,C336V13,C769V13,C1122V13,V13C336,V13C769,V13C1122,SI13,end_vn13);
V14:VNPU3_3 port map (start_vn,clk,rst,Lc14,C337V14,C770V14,C1123V14,V14C337,V14C770,V14C1123,SI14,end_vn14);
V15:VNPU3_3 port map (start_vn,clk,rst,Lc15,C338V15,C771V15,C1124V15,V15C338,V15C771,V15C1124,SI15,end_vn15);
V16:VNPU3_3 port map (start_vn,clk,rst,Lc16,C339V16,C772V16,C1125V16,V16C339,V16C772,V16C1125,SI16,end_vn16);
V17:VNPU3_3 port map (start_vn,clk,rst,Lc17,C340V17,C773V17,C1126V17,V17C340,V17C773,V17C1126,SI17,end_vn17);
V18:VNPU3_3 port map (start_vn,clk,rst,Lc18,C341V18,C774V18,C1127V18,V18C341,V18C774,V18C1127,SI18,end_vn18);
V19:VNPU3_3 port map (start_vn,clk,rst,Lc19,C342V19,C775V19,C1128V19,V19C342,V19C775,V19C1128,SI19,end_vn19);
V20:VNPU3_3 port map (start_vn,clk,rst,Lc20,C343V20,C776V20,C1129V20,V20C343,V20C776,V20C1129,SI20,end_vn20);
V21:VNPU3_3 port map (start_vn,clk,rst,Lc21,C344V21,C777V21,C1130V21,V21C344,V21C777,V21C1130,SI21,end_vn21);
V22:VNPU3_3 port map (start_vn,clk,rst,Lc22,C345V22,C778V22,C1131V22,V22C345,V22C778,V22C1131,SI22,end_vn22);
V23:VNPU3_3 port map (start_vn,clk,rst,Lc23,C346V23,C779V23,C1132V23,V23C346,V23C779,V23C1132,SI23,end_vn23);
V24:VNPU3_3 port map (start_vn,clk,rst,Lc24,C347V24,C780V24,C1133V24,V24C347,V24C780,V24C1133,SI24,end_vn24);
V25:VNPU3_3 port map (start_vn,clk,rst,Lc25,C348V25,C781V25,C1134V25,V25C348,V25C781,V25C1134,SI25,end_vn25);
V26:VNPU3_3 port map (start_vn,clk,rst,Lc26,C349V26,C782V26,C1135V26,V26C349,V26C782,V26C1135,SI26,end_vn26);
V27:VNPU3_3 port map (start_vn,clk,rst,Lc27,C350V27,C783V27,C1136V27,V27C350,V27C783,V27C1136,SI27,end_vn27);
V28:VNPU3_3 port map (start_vn,clk,rst,Lc28,C351V28,C784V28,C1137V28,V28C351,V28C784,V28C1137,SI28,end_vn28);
V29:VNPU3_3 port map (start_vn,clk,rst,Lc29,C352V29,C785V29,C1138V29,V29C352,V29C785,V29C1138,SI29,end_vn29);
V30:VNPU3_3 port map (start_vn,clk,rst,Lc30,C353V30,C786V30,C1139V30,V30C353,V30C786,V30C1139,SI30,end_vn30);
V31:VNPU3_3 port map (start_vn,clk,rst,Lc31,C354V31,C787V31,C1140V31,V31C354,V31C787,V31C1140,SI31,end_vn31);
V32:VNPU3_3 port map (start_vn,clk,rst,Lc32,C355V32,C788V32,C1141V32,V32C355,V32C788,V32C1141,SI32,end_vn32);
V33:VNPU3_3 port map (start_vn,clk,rst,Lc33,C356V33,C789V33,C1142V33,V33C356,V33C789,V33C1142,SI33,end_vn33);
V34:VNPU3_3 port map (start_vn,clk,rst,Lc34,C357V34,C790V34,C1143V34,V34C357,V34C790,V34C1143,SI34,end_vn34);
V35:VNPU3_3 port map (start_vn,clk,rst,Lc35,C358V35,C791V35,C1144V35,V35C358,V35C791,V35C1144,SI35,end_vn35);
V36:VNPU3_3 port map (start_vn,clk,rst,Lc36,C359V36,C792V36,C1145V36,V36C359,V36C792,V36C1145,SI36,end_vn36);
V37:VNPU3_3 port map (start_vn,clk,rst,Lc37,C360V37,C793V37,C1146V37,V37C360,V37C793,V37C1146,SI37,end_vn37);
V38:VNPU3_3 port map (start_vn,clk,rst,Lc38,C361V38,C794V38,C1147V38,V38C361,V38C794,V38C1147,SI38,end_vn38);
V39:VNPU3_3 port map (start_vn,clk,rst,Lc39,C362V39,C795V39,C1148V39,V39C362,V39C795,V39C1148,SI39,end_vn39);
V40:VNPU3_3 port map (start_vn,clk,rst,Lc40,C363V40,C796V40,C1149V40,V40C363,V40C796,V40C1149,SI40,end_vn40);
V41:VNPU3_3 port map (start_vn,clk,rst,Lc41,C364V41,C797V41,C1150V41,V41C364,V41C797,V41C1150,SI41,end_vn41);
V42:VNPU3_3 port map (start_vn,clk,rst,Lc42,C365V42,C798V42,C1151V42,V42C365,V42C798,V42C1151,SI42,end_vn42);
V43:VNPU3_3 port map (start_vn,clk,rst,Lc43,C366V43,C799V43,C1152V43,V43C366,V43C799,V43C1152,SI43,end_vn43);
V44:VNPU3_3 port map (start_vn,clk,rst,Lc44,C367V44,C800V44,C1057V44,V44C367,V44C800,V44C1057,SI44,end_vn44);
V45:VNPU3_3 port map (start_vn,clk,rst,Lc45,C368V45,C801V45,C1058V45,V45C368,V45C801,V45C1058,SI45,end_vn45);
V46:VNPU3_3 port map (start_vn,clk,rst,Lc46,C369V46,C802V46,C1059V46,V46C369,V46C802,V46C1059,SI46,end_vn46);
V47:VNPU3_3 port map (start_vn,clk,rst,Lc47,C370V47,C803V47,C1060V47,V47C370,V47C803,V47C1060,SI47,end_vn47);
V48:VNPU3_3 port map (start_vn,clk,rst,Lc48,C371V48,C804V48,C1061V48,V48C371,V48C804,V48C1061,SI48,end_vn48);
V49:VNPU3_3 port map (start_vn,clk,rst,Lc49,C372V49,C805V49,C1062V49,V49C372,V49C805,V49C1062,SI49,end_vn49);
V50:VNPU3_3 port map (start_vn,clk,rst,Lc50,C373V50,C806V50,C1063V50,V50C373,V50C806,V50C1063,SI50,end_vn50);
V51:VNPU3_3 port map (start_vn,clk,rst,Lc51,C374V51,C807V51,C1064V51,V51C374,V51C807,V51C1064,SI51,end_vn51);
V52:VNPU3_3 port map (start_vn,clk,rst,Lc52,C375V52,C808V52,C1065V52,V52C375,V52C808,V52C1065,SI52,end_vn52);
V53:VNPU3_3 port map (start_vn,clk,rst,Lc53,C376V53,C809V53,C1066V53,V53C376,V53C809,V53C1066,SI53,end_vn53);
V54:VNPU3_3 port map (start_vn,clk,rst,Lc54,C377V54,C810V54,C1067V54,V54C377,V54C810,V54C1067,SI54,end_vn54);
V55:VNPU3_3 port map (start_vn,clk,rst,Lc55,C378V55,C811V55,C1068V55,V55C378,V55C811,V55C1068,SI55,end_vn55);
V56:VNPU3_3 port map (start_vn,clk,rst,Lc56,C379V56,C812V56,C1069V56,V56C379,V56C812,V56C1069,SI56,end_vn56);
V57:VNPU3_3 port map (start_vn,clk,rst,Lc57,C380V57,C813V57,C1070V57,V57C380,V57C813,V57C1070,SI57,end_vn57);
V58:VNPU3_3 port map (start_vn,clk,rst,Lc58,C381V58,C814V58,C1071V58,V58C381,V58C814,V58C1071,SI58,end_vn58);
V59:VNPU3_3 port map (start_vn,clk,rst,Lc59,C382V59,C815V59,C1072V59,V59C382,V59C815,V59C1072,SI59,end_vn59);
V60:VNPU3_3 port map (start_vn,clk,rst,Lc60,C383V60,C816V60,C1073V60,V60C383,V60C816,V60C1073,SI60,end_vn60);
V61:VNPU3_3 port map (start_vn,clk,rst,Lc61,C384V61,C817V61,C1074V61,V61C384,V61C817,V61C1074,SI61,end_vn61);
V62:VNPU3_3 port map (start_vn,clk,rst,Lc62,C289V62,C818V62,C1075V62,V62C289,V62C818,V62C1075,SI62,end_vn62);
V63:VNPU3_3 port map (start_vn,clk,rst,Lc63,C290V63,C819V63,C1076V63,V63C290,V63C819,V63C1076,SI63,end_vn63);
V64:VNPU3_3 port map (start_vn,clk,rst,Lc64,C291V64,C820V64,C1077V64,V64C291,V64C820,V64C1077,SI64,end_vn64);
V65:VNPU3_3 port map (start_vn,clk,rst,Lc65,C292V65,C821V65,C1078V65,V65C292,V65C821,V65C1078,SI65,end_vn65);
V66:VNPU3_3 port map (start_vn,clk,rst,Lc66,C293V66,C822V66,C1079V66,V66C293,V66C822,V66C1079,SI66,end_vn66);
V67:VNPU3_3 port map (start_vn,clk,rst,Lc67,C294V67,C823V67,C1080V67,V67C294,V67C823,V67C1080,SI67,end_vn67);
V68:VNPU3_3 port map (start_vn,clk,rst,Lc68,C295V68,C824V68,C1081V68,V68C295,V68C824,V68C1081,SI68,end_vn68);
V69:VNPU3_3 port map (start_vn,clk,rst,Lc69,C296V69,C825V69,C1082V69,V69C296,V69C825,V69C1082,SI69,end_vn69);
V70:VNPU3_3 port map (start_vn,clk,rst,Lc70,C297V70,C826V70,C1083V70,V70C297,V70C826,V70C1083,SI70,end_vn70);
V71:VNPU3_3 port map (start_vn,clk,rst,Lc71,C298V71,C827V71,C1084V71,V71C298,V71C827,V71C1084,SI71,end_vn71);
V72:VNPU3_3 port map (start_vn,clk,rst,Lc72,C299V72,C828V72,C1085V72,V72C299,V72C828,V72C1085,SI72,end_vn72);
V73:VNPU3_3 port map (start_vn,clk,rst,Lc73,C300V73,C829V73,C1086V73,V73C300,V73C829,V73C1086,SI73,end_vn73);
V74:VNPU3_3 port map (start_vn,clk,rst,Lc74,C301V74,C830V74,C1087V74,V74C301,V74C830,V74C1087,SI74,end_vn74);
V75:VNPU3_3 port map (start_vn,clk,rst,Lc75,C302V75,C831V75,C1088V75,V75C302,V75C831,V75C1088,SI75,end_vn75);
V76:VNPU3_3 port map (start_vn,clk,rst,Lc76,C303V76,C832V76,C1089V76,V76C303,V76C832,V76C1089,SI76,end_vn76);
V77:VNPU3_3 port map (start_vn,clk,rst,Lc77,C304V77,C833V77,C1090V77,V77C304,V77C833,V77C1090,SI77,end_vn77);
V78:VNPU3_3 port map (start_vn,clk,rst,Lc78,C305V78,C834V78,C1091V78,V78C305,V78C834,V78C1091,SI78,end_vn78);
V79:VNPU3_3 port map (start_vn,clk,rst,Lc79,C306V79,C835V79,C1092V79,V79C306,V79C835,V79C1092,SI79,end_vn79);
V80:VNPU3_3 port map (start_vn,clk,rst,Lc80,C307V80,C836V80,C1093V80,V80C307,V80C836,V80C1093,SI80,end_vn80);
V81:VNPU3_3 port map (start_vn,clk,rst,Lc81,C308V81,C837V81,C1094V81,V81C308,V81C837,V81C1094,SI81,end_vn81);
V82:VNPU3_3 port map (start_vn,clk,rst,Lc82,C309V82,C838V82,C1095V82,V82C309,V82C838,V82C1095,SI82,end_vn82);
V83:VNPU3_3 port map (start_vn,clk,rst,Lc83,C310V83,C839V83,C1096V83,V83C310,V83C839,V83C1096,SI83,end_vn83);
V84:VNPU3_3 port map (start_vn,clk,rst,Lc84,C311V84,C840V84,C1097V84,V84C311,V84C840,V84C1097,SI84,end_vn84);
V85:VNPU3_3 port map (start_vn,clk,rst,Lc85,C312V85,C841V85,C1098V85,V85C312,V85C841,V85C1098,SI85,end_vn85);
V86:VNPU3_3 port map (start_vn,clk,rst,Lc86,C313V86,C842V86,C1099V86,V86C313,V86C842,V86C1099,SI86,end_vn86);
V87:VNPU3_3 port map (start_vn,clk,rst,Lc87,C314V87,C843V87,C1100V87,V87C314,V87C843,V87C1100,SI87,end_vn87);
V88:VNPU3_3 port map (start_vn,clk,rst,Lc88,C315V88,C844V88,C1101V88,V88C315,V88C844,V88C1101,SI88,end_vn88);
V89:VNPU3_3 port map (start_vn,clk,rst,Lc89,C316V89,C845V89,C1102V89,V89C316,V89C845,V89C1102,SI89,end_vn89);
V90:VNPU3_3 port map (start_vn,clk,rst,Lc90,C317V90,C846V90,C1103V90,V90C317,V90C846,V90C1103,SI90,end_vn90);
V91:VNPU3_3 port map (start_vn,clk,rst,Lc91,C318V91,C847V91,C1104V91,V91C318,V91C847,V91C1104,SI91,end_vn91);
V92:VNPU3_3 port map (start_vn,clk,rst,Lc92,C319V92,C848V92,C1105V92,V92C319,V92C848,V92C1105,SI92,end_vn92);
V93:VNPU3_3 port map (start_vn,clk,rst,Lc93,C320V93,C849V93,C1106V93,V93C320,V93C849,V93C1106,SI93,end_vn93);
V94:VNPU3_3 port map (start_vn,clk,rst,Lc94,C321V94,C850V94,C1107V94,V94C321,V94C850,V94C1107,SI94,end_vn94);
V95:VNPU3_3 port map (start_vn,clk,rst,Lc95,C322V95,C851V95,C1108V95,V95C322,V95C851,V95C1108,SI95,end_vn95);
V96:VNPU3_3 port map (start_vn,clk,rst,Lc96,C323V96,C852V96,C1109V96,V96C323,V96C852,V96C1109,SI96,end_vn96);
V97:VNPU3_3 port map (start_vn,clk,rst,Lc97,C3V97,C166V97,C758V97,V97C3,V97C166,V97C758,SI97,end_vn97);
V98:VNPU3_3 port map (start_vn,clk,rst,Lc98,C4V98,C167V98,C759V98,V98C4,V98C167,V98C759,SI98,end_vn98);
V99:VNPU3_3 port map (start_vn,clk,rst,Lc99,C5V99,C168V99,C760V99,V99C5,V99C168,V99C760,SI99,end_vn99);
V100:VNPU3_3 port map (start_vn,clk,rst,Lc100,C6V100,C169V100,C761V100,V100C6,V100C169,V100C761,SI100,end_vn100);
V101:VNPU3_3 port map (start_vn,clk,rst,Lc101,C7V101,C170V101,C762V101,V101C7,V101C170,V101C762,SI101,end_vn101);
V102:VNPU3_3 port map (start_vn,clk,rst,Lc102,C8V102,C171V102,C763V102,V102C8,V102C171,V102C763,SI102,end_vn102);
V103:VNPU3_3 port map (start_vn,clk,rst,Lc103,C9V103,C172V103,C764V103,V103C9,V103C172,V103C764,SI103,end_vn103);
V104:VNPU3_3 port map (start_vn,clk,rst,Lc104,C10V104,C173V104,C765V104,V104C10,V104C173,V104C765,SI104,end_vn104);
V105:VNPU3_3 port map (start_vn,clk,rst,Lc105,C11V105,C174V105,C766V105,V105C11,V105C174,V105C766,SI105,end_vn105);
V106:VNPU3_3 port map (start_vn,clk,rst,Lc106,C12V106,C175V106,C767V106,V106C12,V106C175,V106C767,SI106,end_vn106);
V107:VNPU3_3 port map (start_vn,clk,rst,Lc107,C13V107,C176V107,C768V107,V107C13,V107C176,V107C768,SI107,end_vn107);
V108:VNPU3_3 port map (start_vn,clk,rst,Lc108,C14V108,C177V108,C673V108,V108C14,V108C177,V108C673,SI108,end_vn108);
V109:VNPU3_3 port map (start_vn,clk,rst,Lc109,C15V109,C178V109,C674V109,V109C15,V109C178,V109C674,SI109,end_vn109);
V110:VNPU3_3 port map (start_vn,clk,rst,Lc110,C16V110,C179V110,C675V110,V110C16,V110C179,V110C675,SI110,end_vn110);
V111:VNPU3_3 port map (start_vn,clk,rst,Lc111,C17V111,C180V111,C676V111,V111C17,V111C180,V111C676,SI111,end_vn111);
V112:VNPU3_3 port map (start_vn,clk,rst,Lc112,C18V112,C181V112,C677V112,V112C18,V112C181,V112C677,SI112,end_vn112);
V113:VNPU3_3 port map (start_vn,clk,rst,Lc113,C19V113,C182V113,C678V113,V113C19,V113C182,V113C678,SI113,end_vn113);
V114:VNPU3_3 port map (start_vn,clk,rst,Lc114,C20V114,C183V114,C679V114,V114C20,V114C183,V114C679,SI114,end_vn114);
V115:VNPU3_3 port map (start_vn,clk,rst,Lc115,C21V115,C184V115,C680V115,V115C21,V115C184,V115C680,SI115,end_vn115);
V116:VNPU3_3 port map (start_vn,clk,rst,Lc116,C22V116,C185V116,C681V116,V116C22,V116C185,V116C681,SI116,end_vn116);
V117:VNPU3_3 port map (start_vn,clk,rst,Lc117,C23V117,C186V117,C682V117,V117C23,V117C186,V117C682,SI117,end_vn117);
V118:VNPU3_3 port map (start_vn,clk,rst,Lc118,C24V118,C187V118,C683V118,V118C24,V118C187,V118C683,SI118,end_vn118);
V119:VNPU3_3 port map (start_vn,clk,rst,Lc119,C25V119,C188V119,C684V119,V119C25,V119C188,V119C684,SI119,end_vn119);
V120:VNPU3_3 port map (start_vn,clk,rst,Lc120,C26V120,C189V120,C685V120,V120C26,V120C189,V120C685,SI120,end_vn120);
V121:VNPU3_3 port map (start_vn,clk,rst,Lc121,C27V121,C190V121,C686V121,V121C27,V121C190,V121C686,SI121,end_vn121);
V122:VNPU3_3 port map (start_vn,clk,rst,Lc122,C28V122,C191V122,C687V122,V122C28,V122C191,V122C687,SI122,end_vn122);
V123:VNPU3_3 port map (start_vn,clk,rst,Lc123,C29V123,C192V123,C688V123,V123C29,V123C192,V123C688,SI123,end_vn123);
V124:VNPU3_3 port map (start_vn,clk,rst,Lc124,C30V124,C97V124,C689V124,V124C30,V124C97,V124C689,SI124,end_vn124);
V125:VNPU3_3 port map (start_vn,clk,rst,Lc125,C31V125,C98V125,C690V125,V125C31,V125C98,V125C690,SI125,end_vn125);
V126:VNPU3_3 port map (start_vn,clk,rst,Lc126,C32V126,C99V126,C691V126,V126C32,V126C99,V126C691,SI126,end_vn126);
V127:VNPU3_3 port map (start_vn,clk,rst,Lc127,C33V127,C100V127,C692V127,V127C33,V127C100,V127C692,SI127,end_vn127);
V128:VNPU3_3 port map (start_vn,clk,rst,Lc128,C34V128,C101V128,C693V128,V128C34,V128C101,V128C693,SI128,end_vn128);
V129:VNPU3_3 port map (start_vn,clk,rst,Lc129,C35V129,C102V129,C694V129,V129C35,V129C102,V129C694,SI129,end_vn129);
V130:VNPU3_3 port map (start_vn,clk,rst,Lc130,C36V130,C103V130,C695V130,V130C36,V130C103,V130C695,SI130,end_vn130);
V131:VNPU3_3 port map (start_vn,clk,rst,Lc131,C37V131,C104V131,C696V131,V131C37,V131C104,V131C696,SI131,end_vn131);
V132:VNPU3_3 port map (start_vn,clk,rst,Lc132,C38V132,C105V132,C697V132,V132C38,V132C105,V132C697,SI132,end_vn132);
V133:VNPU3_3 port map (start_vn,clk,rst,Lc133,C39V133,C106V133,C698V133,V133C39,V133C106,V133C698,SI133,end_vn133);
V134:VNPU3_3 port map (start_vn,clk,rst,Lc134,C40V134,C107V134,C699V134,V134C40,V134C107,V134C699,SI134,end_vn134);
V135:VNPU3_3 port map (start_vn,clk,rst,Lc135,C41V135,C108V135,C700V135,V135C41,V135C108,V135C700,SI135,end_vn135);
V136:VNPU3_3 port map (start_vn,clk,rst,Lc136,C42V136,C109V136,C701V136,V136C42,V136C109,V136C701,SI136,end_vn136);
V137:VNPU3_3 port map (start_vn,clk,rst,Lc137,C43V137,C110V137,C702V137,V137C43,V137C110,V137C702,SI137,end_vn137);
V138:VNPU3_3 port map (start_vn,clk,rst,Lc138,C44V138,C111V138,C703V138,V138C44,V138C111,V138C703,SI138,end_vn138);
V139:VNPU3_3 port map (start_vn,clk,rst,Lc139,C45V139,C112V139,C704V139,V139C45,V139C112,V139C704,SI139,end_vn139);
V140:VNPU3_3 port map (start_vn,clk,rst,Lc140,C46V140,C113V140,C705V140,V140C46,V140C113,V140C705,SI140,end_vn140);
V141:VNPU3_3 port map (start_vn,clk,rst,Lc141,C47V141,C114V141,C706V141,V141C47,V141C114,V141C706,SI141,end_vn141);
V142:VNPU3_3 port map (start_vn,clk,rst,Lc142,C48V142,C115V142,C707V142,V142C48,V142C115,V142C707,SI142,end_vn142);
V143:VNPU3_3 port map (start_vn,clk,rst,Lc143,C49V143,C116V143,C708V143,V143C49,V143C116,V143C708,SI143,end_vn143);
V144:VNPU3_3 port map (start_vn,clk,rst,Lc144,C50V144,C117V144,C709V144,V144C50,V144C117,V144C709,SI144,end_vn144);
V145:VNPU3_3 port map (start_vn,clk,rst,Lc145,C51V145,C118V145,C710V145,V145C51,V145C118,V145C710,SI145,end_vn145);
V146:VNPU3_3 port map (start_vn,clk,rst,Lc146,C52V146,C119V146,C711V146,V146C52,V146C119,V146C711,SI146,end_vn146);
V147:VNPU3_3 port map (start_vn,clk,rst,Lc147,C53V147,C120V147,C712V147,V147C53,V147C120,V147C712,SI147,end_vn147);
V148:VNPU3_3 port map (start_vn,clk,rst,Lc148,C54V148,C121V148,C713V148,V148C54,V148C121,V148C713,SI148,end_vn148);
V149:VNPU3_3 port map (start_vn,clk,rst,Lc149,C55V149,C122V149,C714V149,V149C55,V149C122,V149C714,SI149,end_vn149);
V150:VNPU3_3 port map (start_vn,clk,rst,Lc150,C56V150,C123V150,C715V150,V150C56,V150C123,V150C715,SI150,end_vn150);
V151:VNPU3_3 port map (start_vn,clk,rst,Lc151,C57V151,C124V151,C716V151,V151C57,V151C124,V151C716,SI151,end_vn151);
V152:VNPU3_3 port map (start_vn,clk,rst,Lc152,C58V152,C125V152,C717V152,V152C58,V152C125,V152C717,SI152,end_vn152);
V153:VNPU3_3 port map (start_vn,clk,rst,Lc153,C59V153,C126V153,C718V153,V153C59,V153C126,V153C718,SI153,end_vn153);
V154:VNPU3_3 port map (start_vn,clk,rst,Lc154,C60V154,C127V154,C719V154,V154C60,V154C127,V154C719,SI154,end_vn154);
V155:VNPU3_3 port map (start_vn,clk,rst,Lc155,C61V155,C128V155,C720V155,V155C61,V155C128,V155C720,SI155,end_vn155);
V156:VNPU3_3 port map (start_vn,clk,rst,Lc156,C62V156,C129V156,C721V156,V156C62,V156C129,V156C721,SI156,end_vn156);
V157:VNPU3_3 port map (start_vn,clk,rst,Lc157,C63V157,C130V157,C722V157,V157C63,V157C130,V157C722,SI157,end_vn157);
V158:VNPU3_3 port map (start_vn,clk,rst,Lc158,C64V158,C131V158,C723V158,V158C64,V158C131,V158C723,SI158,end_vn158);
V159:VNPU3_3 port map (start_vn,clk,rst,Lc159,C65V159,C132V159,C724V159,V159C65,V159C132,V159C724,SI159,end_vn159);
V160:VNPU3_3 port map (start_vn,clk,rst,Lc160,C66V160,C133V160,C725V160,V160C66,V160C133,V160C725,SI160,end_vn160);
V161:VNPU3_3 port map (start_vn,clk,rst,Lc161,C67V161,C134V161,C726V161,V161C67,V161C134,V161C726,SI161,end_vn161);
V162:VNPU3_3 port map (start_vn,clk,rst,Lc162,C68V162,C135V162,C727V162,V162C68,V162C135,V162C727,SI162,end_vn162);
V163:VNPU3_3 port map (start_vn,clk,rst,Lc163,C69V163,C136V163,C728V163,V163C69,V163C136,V163C728,SI163,end_vn163);
V164:VNPU3_3 port map (start_vn,clk,rst,Lc164,C70V164,C137V164,C729V164,V164C70,V164C137,V164C729,SI164,end_vn164);
V165:VNPU3_3 port map (start_vn,clk,rst,Lc165,C71V165,C138V165,C730V165,V165C71,V165C138,V165C730,SI165,end_vn165);
V166:VNPU3_3 port map (start_vn,clk,rst,Lc166,C72V166,C139V166,C731V166,V166C72,V166C139,V166C731,SI166,end_vn166);
V167:VNPU3_3 port map (start_vn,clk,rst,Lc167,C73V167,C140V167,C732V167,V167C73,V167C140,V167C732,SI167,end_vn167);
V168:VNPU3_3 port map (start_vn,clk,rst,Lc168,C74V168,C141V168,C733V168,V168C74,V168C141,V168C733,SI168,end_vn168);
V169:VNPU3_3 port map (start_vn,clk,rst,Lc169,C75V169,C142V169,C734V169,V169C75,V169C142,V169C734,SI169,end_vn169);
V170:VNPU3_3 port map (start_vn,clk,rst,Lc170,C76V170,C143V170,C735V170,V170C76,V170C143,V170C735,SI170,end_vn170);
V171:VNPU3_3 port map (start_vn,clk,rst,Lc171,C77V171,C144V171,C736V171,V171C77,V171C144,V171C736,SI171,end_vn171);
V172:VNPU3_3 port map (start_vn,clk,rst,Lc172,C78V172,C145V172,C737V172,V172C78,V172C145,V172C737,SI172,end_vn172);
V173:VNPU3_3 port map (start_vn,clk,rst,Lc173,C79V173,C146V173,C738V173,V173C79,V173C146,V173C738,SI173,end_vn173);
V174:VNPU3_3 port map (start_vn,clk,rst,Lc174,C80V174,C147V174,C739V174,V174C80,V174C147,V174C739,SI174,end_vn174);
V175:VNPU3_3 port map (start_vn,clk,rst,Lc175,C81V175,C148V175,C740V175,V175C81,V175C148,V175C740,SI175,end_vn175);
V176:VNPU3_3 port map (start_vn,clk,rst,Lc176,C82V176,C149V176,C741V176,V176C82,V176C149,V176C741,SI176,end_vn176);
V177:VNPU3_3 port map (start_vn,clk,rst,Lc177,C83V177,C150V177,C742V177,V177C83,V177C150,V177C742,SI177,end_vn177);
V178:VNPU3_3 port map (start_vn,clk,rst,Lc178,C84V178,C151V178,C743V178,V178C84,V178C151,V178C743,SI178,end_vn178);
V179:VNPU3_3 port map (start_vn,clk,rst,Lc179,C85V179,C152V179,C744V179,V179C85,V179C152,V179C744,SI179,end_vn179);
V180:VNPU3_3 port map (start_vn,clk,rst,Lc180,C86V180,C153V180,C745V180,V180C86,V180C153,V180C745,SI180,end_vn180);
V181:VNPU3_3 port map (start_vn,clk,rst,Lc181,C87V181,C154V181,C746V181,V181C87,V181C154,V181C746,SI181,end_vn181);
V182:VNPU3_3 port map (start_vn,clk,rst,Lc182,C88V182,C155V182,C747V182,V182C88,V182C155,V182C747,SI182,end_vn182);
V183:VNPU3_3 port map (start_vn,clk,rst,Lc183,C89V183,C156V183,C748V183,V183C89,V183C156,V183C748,SI183,end_vn183);
V184:VNPU3_3 port map (start_vn,clk,rst,Lc184,C90V184,C157V184,C749V184,V184C90,V184C157,V184C749,SI184,end_vn184);
V185:VNPU3_3 port map (start_vn,clk,rst,Lc185,C91V185,C158V185,C750V185,V185C91,V185C158,V185C750,SI185,end_vn185);
V186:VNPU3_3 port map (start_vn,clk,rst,Lc186,C92V186,C159V186,C751V186,V186C92,V186C159,V186C751,SI186,end_vn186);
V187:VNPU3_3 port map (start_vn,clk,rst,Lc187,C93V187,C160V187,C752V187,V187C93,V187C160,V187C752,SI187,end_vn187);
V188:VNPU3_3 port map (start_vn,clk,rst,Lc188,C94V188,C161V188,C753V188,V188C94,V188C161,V188C753,SI188,end_vn188);
V189:VNPU3_3 port map (start_vn,clk,rst,Lc189,C95V189,C162V189,C754V189,V189C95,V189C162,V189C754,SI189,end_vn189);
V190:VNPU3_3 port map (start_vn,clk,rst,Lc190,C96V190,C163V190,C755V190,V190C96,V190C163,V190C755,SI190,end_vn190);
V191:VNPU3_3 port map (start_vn,clk,rst,Lc191,C1V191,C164V191,C756V191,V191C1,V191C164,V191C756,SI191,end_vn191);
V192:VNPU3_3 port map (start_vn,clk,rst,Lc192,C2V192,C165V192,C757V192,V192C2,V192C165,V192C757,SI192,end_vn192);
V193:VNPU6_6 port map (start_vn,clk,rst,Lc193,C24V193,C338V193,C442V193,C578V193,C696V193,C1050V193,V193C24,V193C338,V193C442,V193C578,V193C696,V193C1050,SI193,end_vn193);
V194:VNPU6_6 port map (start_vn,clk,rst,Lc194,C25V194,C339V194,C443V194,C579V194,C697V194,C1051V194,V194C25,V194C339,V194C443,V194C579,V194C697,V194C1051,SI194,end_vn194);
V195:VNPU6_6 port map (start_vn,clk,rst,Lc195,C26V195,C340V195,C444V195,C580V195,C698V195,C1052V195,V195C26,V195C340,V195C444,V195C580,V195C698,V195C1052,SI195,end_vn195);
V196:VNPU6_6 port map (start_vn,clk,rst,Lc196,C27V196,C341V196,C445V196,C581V196,C699V196,C1053V196,V196C27,V196C341,V196C445,V196C581,V196C699,V196C1053,SI196,end_vn196);
V197:VNPU6_6 port map (start_vn,clk,rst,Lc197,C28V197,C342V197,C446V197,C582V197,C700V197,C1054V197,V197C28,V197C342,V197C446,V197C582,V197C700,V197C1054,SI197,end_vn197);
V198:VNPU6_6 port map (start_vn,clk,rst,Lc198,C29V198,C343V198,C447V198,C583V198,C701V198,C1055V198,V198C29,V198C343,V198C447,V198C583,V198C701,V198C1055,SI198,end_vn198);
V199:VNPU6_6 port map (start_vn,clk,rst,Lc199,C30V199,C344V199,C448V199,C584V199,C702V199,C1056V199,V199C30,V199C344,V199C448,V199C584,V199C702,V199C1056,SI199,end_vn199);
V200:VNPU6_6 port map (start_vn,clk,rst,Lc200,C31V200,C345V200,C449V200,C585V200,C703V200,C961V200,V200C31,V200C345,V200C449,V200C585,V200C703,V200C961,SI200,end_vn200);
V201:VNPU6_6 port map (start_vn,clk,rst,Lc201,C32V201,C346V201,C450V201,C586V201,C704V201,C962V201,V201C32,V201C346,V201C450,V201C586,V201C704,V201C962,SI201,end_vn201);
V202:VNPU6_6 port map (start_vn,clk,rst,Lc202,C33V202,C347V202,C451V202,C587V202,C705V202,C963V202,V202C33,V202C347,V202C451,V202C587,V202C705,V202C963,SI202,end_vn202);
V203:VNPU6_6 port map (start_vn,clk,rst,Lc203,C34V203,C348V203,C452V203,C588V203,C706V203,C964V203,V203C34,V203C348,V203C452,V203C588,V203C706,V203C964,SI203,end_vn203);
V204:VNPU6_6 port map (start_vn,clk,rst,Lc204,C35V204,C349V204,C453V204,C589V204,C707V204,C965V204,V204C35,V204C349,V204C453,V204C589,V204C707,V204C965,SI204,end_vn204);
V205:VNPU6_6 port map (start_vn,clk,rst,Lc205,C36V205,C350V205,C454V205,C590V205,C708V205,C966V205,V205C36,V205C350,V205C454,V205C590,V205C708,V205C966,SI205,end_vn205);
V206:VNPU6_6 port map (start_vn,clk,rst,Lc206,C37V206,C351V206,C455V206,C591V206,C709V206,C967V206,V206C37,V206C351,V206C455,V206C591,V206C709,V206C967,SI206,end_vn206);
V207:VNPU6_6 port map (start_vn,clk,rst,Lc207,C38V207,C352V207,C456V207,C592V207,C710V207,C968V207,V207C38,V207C352,V207C456,V207C592,V207C710,V207C968,SI207,end_vn207);
V208:VNPU6_6 port map (start_vn,clk,rst,Lc208,C39V208,C353V208,C457V208,C593V208,C711V208,C969V208,V208C39,V208C353,V208C457,V208C593,V208C711,V208C969,SI208,end_vn208);
V209:VNPU6_6 port map (start_vn,clk,rst,Lc209,C40V209,C354V209,C458V209,C594V209,C712V209,C970V209,V209C40,V209C354,V209C458,V209C594,V209C712,V209C970,SI209,end_vn209);
V210:VNPU6_6 port map (start_vn,clk,rst,Lc210,C41V210,C355V210,C459V210,C595V210,C713V210,C971V210,V210C41,V210C355,V210C459,V210C595,V210C713,V210C971,SI210,end_vn210);
V211:VNPU6_6 port map (start_vn,clk,rst,Lc211,C42V211,C356V211,C460V211,C596V211,C714V211,C972V211,V211C42,V211C356,V211C460,V211C596,V211C714,V211C972,SI211,end_vn211);
V212:VNPU6_6 port map (start_vn,clk,rst,Lc212,C43V212,C357V212,C461V212,C597V212,C715V212,C973V212,V212C43,V212C357,V212C461,V212C597,V212C715,V212C973,SI212,end_vn212);
V213:VNPU6_6 port map (start_vn,clk,rst,Lc213,C44V213,C358V213,C462V213,C598V213,C716V213,C974V213,V213C44,V213C358,V213C462,V213C598,V213C716,V213C974,SI213,end_vn213);
V214:VNPU6_6 port map (start_vn,clk,rst,Lc214,C45V214,C359V214,C463V214,C599V214,C717V214,C975V214,V214C45,V214C359,V214C463,V214C599,V214C717,V214C975,SI214,end_vn214);
V215:VNPU6_6 port map (start_vn,clk,rst,Lc215,C46V215,C360V215,C464V215,C600V215,C718V215,C976V215,V215C46,V215C360,V215C464,V215C600,V215C718,V215C976,SI215,end_vn215);
V216:VNPU6_6 port map (start_vn,clk,rst,Lc216,C47V216,C361V216,C465V216,C601V216,C719V216,C977V216,V216C47,V216C361,V216C465,V216C601,V216C719,V216C977,SI216,end_vn216);
V217:VNPU6_6 port map (start_vn,clk,rst,Lc217,C48V217,C362V217,C466V217,C602V217,C720V217,C978V217,V217C48,V217C362,V217C466,V217C602,V217C720,V217C978,SI217,end_vn217);
V218:VNPU6_6 port map (start_vn,clk,rst,Lc218,C49V218,C363V218,C467V218,C603V218,C721V218,C979V218,V218C49,V218C363,V218C467,V218C603,V218C721,V218C979,SI218,end_vn218);
V219:VNPU6_6 port map (start_vn,clk,rst,Lc219,C50V219,C364V219,C468V219,C604V219,C722V219,C980V219,V219C50,V219C364,V219C468,V219C604,V219C722,V219C980,SI219,end_vn219);
V220:VNPU6_6 port map (start_vn,clk,rst,Lc220,C51V220,C365V220,C469V220,C605V220,C723V220,C981V220,V220C51,V220C365,V220C469,V220C605,V220C723,V220C981,SI220,end_vn220);
V221:VNPU6_6 port map (start_vn,clk,rst,Lc221,C52V221,C366V221,C470V221,C606V221,C724V221,C982V221,V221C52,V221C366,V221C470,V221C606,V221C724,V221C982,SI221,end_vn221);
V222:VNPU6_6 port map (start_vn,clk,rst,Lc222,C53V222,C367V222,C471V222,C607V222,C725V222,C983V222,V222C53,V222C367,V222C471,V222C607,V222C725,V222C983,SI222,end_vn222);
V223:VNPU6_6 port map (start_vn,clk,rst,Lc223,C54V223,C368V223,C472V223,C608V223,C726V223,C984V223,V223C54,V223C368,V223C472,V223C608,V223C726,V223C984,SI223,end_vn223);
V224:VNPU6_6 port map (start_vn,clk,rst,Lc224,C55V224,C369V224,C473V224,C609V224,C727V224,C985V224,V224C55,V224C369,V224C473,V224C609,V224C727,V224C985,SI224,end_vn224);
V225:VNPU6_6 port map (start_vn,clk,rst,Lc225,C56V225,C370V225,C474V225,C610V225,C728V225,C986V225,V225C56,V225C370,V225C474,V225C610,V225C728,V225C986,SI225,end_vn225);
V226:VNPU6_6 port map (start_vn,clk,rst,Lc226,C57V226,C371V226,C475V226,C611V226,C729V226,C987V226,V226C57,V226C371,V226C475,V226C611,V226C729,V226C987,SI226,end_vn226);
V227:VNPU6_6 port map (start_vn,clk,rst,Lc227,C58V227,C372V227,C476V227,C612V227,C730V227,C988V227,V227C58,V227C372,V227C476,V227C612,V227C730,V227C988,SI227,end_vn227);
V228:VNPU6_6 port map (start_vn,clk,rst,Lc228,C59V228,C373V228,C477V228,C613V228,C731V228,C989V228,V228C59,V228C373,V228C477,V228C613,V228C731,V228C989,SI228,end_vn228);
V229:VNPU6_6 port map (start_vn,clk,rst,Lc229,C60V229,C374V229,C478V229,C614V229,C732V229,C990V229,V229C60,V229C374,V229C478,V229C614,V229C732,V229C990,SI229,end_vn229);
V230:VNPU6_6 port map (start_vn,clk,rst,Lc230,C61V230,C375V230,C479V230,C615V230,C733V230,C991V230,V230C61,V230C375,V230C479,V230C615,V230C733,V230C991,SI230,end_vn230);
V231:VNPU6_6 port map (start_vn,clk,rst,Lc231,C62V231,C376V231,C480V231,C616V231,C734V231,C992V231,V231C62,V231C376,V231C480,V231C616,V231C734,V231C992,SI231,end_vn231);
V232:VNPU6_6 port map (start_vn,clk,rst,Lc232,C63V232,C377V232,C385V232,C617V232,C735V232,C993V232,V232C63,V232C377,V232C385,V232C617,V232C735,V232C993,SI232,end_vn232);
V233:VNPU6_6 port map (start_vn,clk,rst,Lc233,C64V233,C378V233,C386V233,C618V233,C736V233,C994V233,V233C64,V233C378,V233C386,V233C618,V233C736,V233C994,SI233,end_vn233);
V234:VNPU6_6 port map (start_vn,clk,rst,Lc234,C65V234,C379V234,C387V234,C619V234,C737V234,C995V234,V234C65,V234C379,V234C387,V234C619,V234C737,V234C995,SI234,end_vn234);
V235:VNPU6_6 port map (start_vn,clk,rst,Lc235,C66V235,C380V235,C388V235,C620V235,C738V235,C996V235,V235C66,V235C380,V235C388,V235C620,V235C738,V235C996,SI235,end_vn235);
V236:VNPU6_6 port map (start_vn,clk,rst,Lc236,C67V236,C381V236,C389V236,C621V236,C739V236,C997V236,V236C67,V236C381,V236C389,V236C621,V236C739,V236C997,SI236,end_vn236);
V237:VNPU6_6 port map (start_vn,clk,rst,Lc237,C68V237,C382V237,C390V237,C622V237,C740V237,C998V237,V237C68,V237C382,V237C390,V237C622,V237C740,V237C998,SI237,end_vn237);
V238:VNPU6_6 port map (start_vn,clk,rst,Lc238,C69V238,C383V238,C391V238,C623V238,C741V238,C999V238,V238C69,V238C383,V238C391,V238C623,V238C741,V238C999,SI238,end_vn238);
V239:VNPU6_6 port map (start_vn,clk,rst,Lc239,C70V239,C384V239,C392V239,C624V239,C742V239,C1000V239,V239C70,V239C384,V239C392,V239C624,V239C742,V239C1000,SI239,end_vn239);
V240:VNPU6_6 port map (start_vn,clk,rst,Lc240,C71V240,C289V240,C393V240,C625V240,C743V240,C1001V240,V240C71,V240C289,V240C393,V240C625,V240C743,V240C1001,SI240,end_vn240);
V241:VNPU6_6 port map (start_vn,clk,rst,Lc241,C72V241,C290V241,C394V241,C626V241,C744V241,C1002V241,V241C72,V241C290,V241C394,V241C626,V241C744,V241C1002,SI241,end_vn241);
V242:VNPU6_6 port map (start_vn,clk,rst,Lc242,C73V242,C291V242,C395V242,C627V242,C745V242,C1003V242,V242C73,V242C291,V242C395,V242C627,V242C745,V242C1003,SI242,end_vn242);
V243:VNPU6_6 port map (start_vn,clk,rst,Lc243,C74V243,C292V243,C396V243,C628V243,C746V243,C1004V243,V243C74,V243C292,V243C396,V243C628,V243C746,V243C1004,SI243,end_vn243);
V244:VNPU6_6 port map (start_vn,clk,rst,Lc244,C75V244,C293V244,C397V244,C629V244,C747V244,C1005V244,V244C75,V244C293,V244C397,V244C629,V244C747,V244C1005,SI244,end_vn244);
V245:VNPU6_6 port map (start_vn,clk,rst,Lc245,C76V245,C294V245,C398V245,C630V245,C748V245,C1006V245,V245C76,V245C294,V245C398,V245C630,V245C748,V245C1006,SI245,end_vn245);
V246:VNPU6_6 port map (start_vn,clk,rst,Lc246,C77V246,C295V246,C399V246,C631V246,C749V246,C1007V246,V246C77,V246C295,V246C399,V246C631,V246C749,V246C1007,SI246,end_vn246);
V247:VNPU6_6 port map (start_vn,clk,rst,Lc247,C78V247,C296V247,C400V247,C632V247,C750V247,C1008V247,V247C78,V247C296,V247C400,V247C632,V247C750,V247C1008,SI247,end_vn247);
V248:VNPU6_6 port map (start_vn,clk,rst,Lc248,C79V248,C297V248,C401V248,C633V248,C751V248,C1009V248,V248C79,V248C297,V248C401,V248C633,V248C751,V248C1009,SI248,end_vn248);
V249:VNPU6_6 port map (start_vn,clk,rst,Lc249,C80V249,C298V249,C402V249,C634V249,C752V249,C1010V249,V249C80,V249C298,V249C402,V249C634,V249C752,V249C1010,SI249,end_vn249);
V250:VNPU6_6 port map (start_vn,clk,rst,Lc250,C81V250,C299V250,C403V250,C635V250,C753V250,C1011V250,V250C81,V250C299,V250C403,V250C635,V250C753,V250C1011,SI250,end_vn250);
V251:VNPU6_6 port map (start_vn,clk,rst,Lc251,C82V251,C300V251,C404V251,C636V251,C754V251,C1012V251,V251C82,V251C300,V251C404,V251C636,V251C754,V251C1012,SI251,end_vn251);
V252:VNPU6_6 port map (start_vn,clk,rst,Lc252,C83V252,C301V252,C405V252,C637V252,C755V252,C1013V252,V252C83,V252C301,V252C405,V252C637,V252C755,V252C1013,SI252,end_vn252);
V253:VNPU6_6 port map (start_vn,clk,rst,Lc253,C84V253,C302V253,C406V253,C638V253,C756V253,C1014V253,V253C84,V253C302,V253C406,V253C638,V253C756,V253C1014,SI253,end_vn253);
V254:VNPU6_6 port map (start_vn,clk,rst,Lc254,C85V254,C303V254,C407V254,C639V254,C757V254,C1015V254,V254C85,V254C303,V254C407,V254C639,V254C757,V254C1015,SI254,end_vn254);
V255:VNPU6_6 port map (start_vn,clk,rst,Lc255,C86V255,C304V255,C408V255,C640V255,C758V255,C1016V255,V255C86,V255C304,V255C408,V255C640,V255C758,V255C1016,SI255,end_vn255);
V256:VNPU6_6 port map (start_vn,clk,rst,Lc256,C87V256,C305V256,C409V256,C641V256,C759V256,C1017V256,V256C87,V256C305,V256C409,V256C641,V256C759,V256C1017,SI256,end_vn256);
V257:VNPU6_6 port map (start_vn,clk,rst,Lc257,C88V257,C306V257,C410V257,C642V257,C760V257,C1018V257,V257C88,V257C306,V257C410,V257C642,V257C760,V257C1018,SI257,end_vn257);
V258:VNPU6_6 port map (start_vn,clk,rst,Lc258,C89V258,C307V258,C411V258,C643V258,C761V258,C1019V258,V258C89,V258C307,V258C411,V258C643,V258C761,V258C1019,SI258,end_vn258);
V259:VNPU6_6 port map (start_vn,clk,rst,Lc259,C90V259,C308V259,C412V259,C644V259,C762V259,C1020V259,V259C90,V259C308,V259C412,V259C644,V259C762,V259C1020,SI259,end_vn259);
V260:VNPU6_6 port map (start_vn,clk,rst,Lc260,C91V260,C309V260,C413V260,C645V260,C763V260,C1021V260,V260C91,V260C309,V260C413,V260C645,V260C763,V260C1021,SI260,end_vn260);
V261:VNPU6_6 port map (start_vn,clk,rst,Lc261,C92V261,C310V261,C414V261,C646V261,C764V261,C1022V261,V261C92,V261C310,V261C414,V261C646,V261C764,V261C1022,SI261,end_vn261);
V262:VNPU6_6 port map (start_vn,clk,rst,Lc262,C93V262,C311V262,C415V262,C647V262,C765V262,C1023V262,V262C93,V262C311,V262C415,V262C647,V262C765,V262C1023,SI262,end_vn262);
V263:VNPU6_6 port map (start_vn,clk,rst,Lc263,C94V263,C312V263,C416V263,C648V263,C766V263,C1024V263,V263C94,V263C312,V263C416,V263C648,V263C766,V263C1024,SI263,end_vn263);
V264:VNPU6_6 port map (start_vn,clk,rst,Lc264,C95V264,C313V264,C417V264,C649V264,C767V264,C1025V264,V264C95,V264C313,V264C417,V264C649,V264C767,V264C1025,SI264,end_vn264);
V265:VNPU6_6 port map (start_vn,clk,rst,Lc265,C96V265,C314V265,C418V265,C650V265,C768V265,C1026V265,V265C96,V265C314,V265C418,V265C650,V265C768,V265C1026,SI265,end_vn265);
V266:VNPU6_6 port map (start_vn,clk,rst,Lc266,C1V266,C315V266,C419V266,C651V266,C673V266,C1027V266,V266C1,V266C315,V266C419,V266C651,V266C673,V266C1027,SI266,end_vn266);
V267:VNPU6_6 port map (start_vn,clk,rst,Lc267,C2V267,C316V267,C420V267,C652V267,C674V267,C1028V267,V267C2,V267C316,V267C420,V267C652,V267C674,V267C1028,SI267,end_vn267);
V268:VNPU6_6 port map (start_vn,clk,rst,Lc268,C3V268,C317V268,C421V268,C653V268,C675V268,C1029V268,V268C3,V268C317,V268C421,V268C653,V268C675,V268C1029,SI268,end_vn268);
V269:VNPU6_6 port map (start_vn,clk,rst,Lc269,C4V269,C318V269,C422V269,C654V269,C676V269,C1030V269,V269C4,V269C318,V269C422,V269C654,V269C676,V269C1030,SI269,end_vn269);
V270:VNPU6_6 port map (start_vn,clk,rst,Lc270,C5V270,C319V270,C423V270,C655V270,C677V270,C1031V270,V270C5,V270C319,V270C423,V270C655,V270C677,V270C1031,SI270,end_vn270);
V271:VNPU6_6 port map (start_vn,clk,rst,Lc271,C6V271,C320V271,C424V271,C656V271,C678V271,C1032V271,V271C6,V271C320,V271C424,V271C656,V271C678,V271C1032,SI271,end_vn271);
V272:VNPU6_6 port map (start_vn,clk,rst,Lc272,C7V272,C321V272,C425V272,C657V272,C679V272,C1033V272,V272C7,V272C321,V272C425,V272C657,V272C679,V272C1033,SI272,end_vn272);
V273:VNPU6_6 port map (start_vn,clk,rst,Lc273,C8V273,C322V273,C426V273,C658V273,C680V273,C1034V273,V273C8,V273C322,V273C426,V273C658,V273C680,V273C1034,SI273,end_vn273);
V274:VNPU6_6 port map (start_vn,clk,rst,Lc274,C9V274,C323V274,C427V274,C659V274,C681V274,C1035V274,V274C9,V274C323,V274C427,V274C659,V274C681,V274C1035,SI274,end_vn274);
V275:VNPU6_6 port map (start_vn,clk,rst,Lc275,C10V275,C324V275,C428V275,C660V275,C682V275,C1036V275,V275C10,V275C324,V275C428,V275C660,V275C682,V275C1036,SI275,end_vn275);
V276:VNPU6_6 port map (start_vn,clk,rst,Lc276,C11V276,C325V276,C429V276,C661V276,C683V276,C1037V276,V276C11,V276C325,V276C429,V276C661,V276C683,V276C1037,SI276,end_vn276);
V277:VNPU6_6 port map (start_vn,clk,rst,Lc277,C12V277,C326V277,C430V277,C662V277,C684V277,C1038V277,V277C12,V277C326,V277C430,V277C662,V277C684,V277C1038,SI277,end_vn277);
V278:VNPU6_6 port map (start_vn,clk,rst,Lc278,C13V278,C327V278,C431V278,C663V278,C685V278,C1039V278,V278C13,V278C327,V278C431,V278C663,V278C685,V278C1039,SI278,end_vn278);
V279:VNPU6_6 port map (start_vn,clk,rst,Lc279,C14V279,C328V279,C432V279,C664V279,C686V279,C1040V279,V279C14,V279C328,V279C432,V279C664,V279C686,V279C1040,SI279,end_vn279);
V280:VNPU6_6 port map (start_vn,clk,rst,Lc280,C15V280,C329V280,C433V280,C665V280,C687V280,C1041V280,V280C15,V280C329,V280C433,V280C665,V280C687,V280C1041,SI280,end_vn280);
V281:VNPU6_6 port map (start_vn,clk,rst,Lc281,C16V281,C330V281,C434V281,C666V281,C688V281,C1042V281,V281C16,V281C330,V281C434,V281C666,V281C688,V281C1042,SI281,end_vn281);
V282:VNPU6_6 port map (start_vn,clk,rst,Lc282,C17V282,C331V282,C435V282,C667V282,C689V282,C1043V282,V282C17,V282C331,V282C435,V282C667,V282C689,V282C1043,SI282,end_vn282);
V283:VNPU6_6 port map (start_vn,clk,rst,Lc283,C18V283,C332V283,C436V283,C668V283,C690V283,C1044V283,V283C18,V283C332,V283C436,V283C668,V283C690,V283C1044,SI283,end_vn283);
V284:VNPU6_6 port map (start_vn,clk,rst,Lc284,C19V284,C333V284,C437V284,C669V284,C691V284,C1045V284,V284C19,V284C333,V284C437,V284C669,V284C691,V284C1045,SI284,end_vn284);
V285:VNPU6_6 port map (start_vn,clk,rst,Lc285,C20V285,C334V285,C438V285,C670V285,C692V285,C1046V285,V285C20,V285C334,V285C438,V285C670,V285C692,V285C1046,SI285,end_vn285);
V286:VNPU6_6 port map (start_vn,clk,rst,Lc286,C21V286,C335V286,C439V286,C671V286,C693V286,C1047V286,V286C21,V286C335,V286C439,V286C671,V286C693,V286C1047,SI286,end_vn286);
V287:VNPU6_6 port map (start_vn,clk,rst,Lc287,C22V287,C336V287,C440V287,C672V287,C694V287,C1048V287,V287C22,V287C336,V287C440,V287C672,V287C694,V287C1048,SI287,end_vn287);
V288:VNPU6_6 port map (start_vn,clk,rst,Lc288,C23V288,C337V288,C441V288,C577V288,C695V288,C1049V288,V288C23,V288C337,V288C441,V288C577,V288C695,V288C1049,SI288,end_vn288);
V289:VNPU3_3 port map (start_vn,clk,rst,Lc289,C265V289,C620V289,C992V289,V289C265,V289C620,V289C992,SI289,end_vn289);
V290:VNPU3_3 port map (start_vn,clk,rst,Lc290,C266V290,C621V290,C993V290,V290C266,V290C621,V290C993,SI290,end_vn290);
V291:VNPU3_3 port map (start_vn,clk,rst,Lc291,C267V291,C622V291,C994V291,V291C267,V291C622,V291C994,SI291,end_vn291);
V292:VNPU3_3 port map (start_vn,clk,rst,Lc292,C268V292,C623V292,C995V292,V292C268,V292C623,V292C995,SI292,end_vn292);
V293:VNPU3_3 port map (start_vn,clk,rst,Lc293,C269V293,C624V293,C996V293,V293C269,V293C624,V293C996,SI293,end_vn293);
V294:VNPU3_3 port map (start_vn,clk,rst,Lc294,C270V294,C625V294,C997V294,V294C270,V294C625,V294C997,SI294,end_vn294);
V295:VNPU3_3 port map (start_vn,clk,rst,Lc295,C271V295,C626V295,C998V295,V295C271,V295C626,V295C998,SI295,end_vn295);
V296:VNPU3_3 port map (start_vn,clk,rst,Lc296,C272V296,C627V296,C999V296,V296C272,V296C627,V296C999,SI296,end_vn296);
V297:VNPU3_3 port map (start_vn,clk,rst,Lc297,C273V297,C628V297,C1000V297,V297C273,V297C628,V297C1000,SI297,end_vn297);
V298:VNPU3_3 port map (start_vn,clk,rst,Lc298,C274V298,C629V298,C1001V298,V298C274,V298C629,V298C1001,SI298,end_vn298);
V299:VNPU3_3 port map (start_vn,clk,rst,Lc299,C275V299,C630V299,C1002V299,V299C275,V299C630,V299C1002,SI299,end_vn299);
V300:VNPU3_3 port map (start_vn,clk,rst,Lc300,C276V300,C631V300,C1003V300,V300C276,V300C631,V300C1003,SI300,end_vn300);
V301:VNPU3_3 port map (start_vn,clk,rst,Lc301,C277V301,C632V301,C1004V301,V301C277,V301C632,V301C1004,SI301,end_vn301);
V302:VNPU3_3 port map (start_vn,clk,rst,Lc302,C278V302,C633V302,C1005V302,V302C278,V302C633,V302C1005,SI302,end_vn302);
V303:VNPU3_3 port map (start_vn,clk,rst,Lc303,C279V303,C634V303,C1006V303,V303C279,V303C634,V303C1006,SI303,end_vn303);
V304:VNPU3_3 port map (start_vn,clk,rst,Lc304,C280V304,C635V304,C1007V304,V304C280,V304C635,V304C1007,SI304,end_vn304);
V305:VNPU3_3 port map (start_vn,clk,rst,Lc305,C281V305,C636V305,C1008V305,V305C281,V305C636,V305C1008,SI305,end_vn305);
V306:VNPU3_3 port map (start_vn,clk,rst,Lc306,C282V306,C637V306,C1009V306,V306C282,V306C637,V306C1009,SI306,end_vn306);
V307:VNPU3_3 port map (start_vn,clk,rst,Lc307,C283V307,C638V307,C1010V307,V307C283,V307C638,V307C1010,SI307,end_vn307);
V308:VNPU3_3 port map (start_vn,clk,rst,Lc308,C284V308,C639V308,C1011V308,V308C284,V308C639,V308C1011,SI308,end_vn308);
V309:VNPU3_3 port map (start_vn,clk,rst,Lc309,C285V309,C640V309,C1012V309,V309C285,V309C640,V309C1012,SI309,end_vn309);
V310:VNPU3_3 port map (start_vn,clk,rst,Lc310,C286V310,C641V310,C1013V310,V310C286,V310C641,V310C1013,SI310,end_vn310);
V311:VNPU3_3 port map (start_vn,clk,rst,Lc311,C287V311,C642V311,C1014V311,V311C287,V311C642,V311C1014,SI311,end_vn311);
V312:VNPU3_3 port map (start_vn,clk,rst,Lc312,C288V312,C643V312,C1015V312,V312C288,V312C643,V312C1015,SI312,end_vn312);
V313:VNPU3_3 port map (start_vn,clk,rst,Lc313,C193V313,C644V313,C1016V313,V313C193,V313C644,V313C1016,SI313,end_vn313);
V314:VNPU3_3 port map (start_vn,clk,rst,Lc314,C194V314,C645V314,C1017V314,V314C194,V314C645,V314C1017,SI314,end_vn314);
V315:VNPU3_3 port map (start_vn,clk,rst,Lc315,C195V315,C646V315,C1018V315,V315C195,V315C646,V315C1018,SI315,end_vn315);
V316:VNPU3_3 port map (start_vn,clk,rst,Lc316,C196V316,C647V316,C1019V316,V316C196,V316C647,V316C1019,SI316,end_vn316);
V317:VNPU3_3 port map (start_vn,clk,rst,Lc317,C197V317,C648V317,C1020V317,V317C197,V317C648,V317C1020,SI317,end_vn317);
V318:VNPU3_3 port map (start_vn,clk,rst,Lc318,C198V318,C649V318,C1021V318,V318C198,V318C649,V318C1021,SI318,end_vn318);
V319:VNPU3_3 port map (start_vn,clk,rst,Lc319,C199V319,C650V319,C1022V319,V319C199,V319C650,V319C1022,SI319,end_vn319);
V320:VNPU3_3 port map (start_vn,clk,rst,Lc320,C200V320,C651V320,C1023V320,V320C200,V320C651,V320C1023,SI320,end_vn320);
V321:VNPU3_3 port map (start_vn,clk,rst,Lc321,C201V321,C652V321,C1024V321,V321C201,V321C652,V321C1024,SI321,end_vn321);
V322:VNPU3_3 port map (start_vn,clk,rst,Lc322,C202V322,C653V322,C1025V322,V322C202,V322C653,V322C1025,SI322,end_vn322);
V323:VNPU3_3 port map (start_vn,clk,rst,Lc323,C203V323,C654V323,C1026V323,V323C203,V323C654,V323C1026,SI323,end_vn323);
V324:VNPU3_3 port map (start_vn,clk,rst,Lc324,C204V324,C655V324,C1027V324,V324C204,V324C655,V324C1027,SI324,end_vn324);
V325:VNPU3_3 port map (start_vn,clk,rst,Lc325,C205V325,C656V325,C1028V325,V325C205,V325C656,V325C1028,SI325,end_vn325);
V326:VNPU3_3 port map (start_vn,clk,rst,Lc326,C206V326,C657V326,C1029V326,V326C206,V326C657,V326C1029,SI326,end_vn326);
V327:VNPU3_3 port map (start_vn,clk,rst,Lc327,C207V327,C658V327,C1030V327,V327C207,V327C658,V327C1030,SI327,end_vn327);
V328:VNPU3_3 port map (start_vn,clk,rst,Lc328,C208V328,C659V328,C1031V328,V328C208,V328C659,V328C1031,SI328,end_vn328);
V329:VNPU3_3 port map (start_vn,clk,rst,Lc329,C209V329,C660V329,C1032V329,V329C209,V329C660,V329C1032,SI329,end_vn329);
V330:VNPU3_3 port map (start_vn,clk,rst,Lc330,C210V330,C661V330,C1033V330,V330C210,V330C661,V330C1033,SI330,end_vn330);
V331:VNPU3_3 port map (start_vn,clk,rst,Lc331,C211V331,C662V331,C1034V331,V331C211,V331C662,V331C1034,SI331,end_vn331);
V332:VNPU3_3 port map (start_vn,clk,rst,Lc332,C212V332,C663V332,C1035V332,V332C212,V332C663,V332C1035,SI332,end_vn332);
V333:VNPU3_3 port map (start_vn,clk,rst,Lc333,C213V333,C664V333,C1036V333,V333C213,V333C664,V333C1036,SI333,end_vn333);
V334:VNPU3_3 port map (start_vn,clk,rst,Lc334,C214V334,C665V334,C1037V334,V334C214,V334C665,V334C1037,SI334,end_vn334);
V335:VNPU3_3 port map (start_vn,clk,rst,Lc335,C215V335,C666V335,C1038V335,V335C215,V335C666,V335C1038,SI335,end_vn335);
V336:VNPU3_3 port map (start_vn,clk,rst,Lc336,C216V336,C667V336,C1039V336,V336C216,V336C667,V336C1039,SI336,end_vn336);
V337:VNPU3_3 port map (start_vn,clk,rst,Lc337,C217V337,C668V337,C1040V337,V337C217,V337C668,V337C1040,SI337,end_vn337);
V338:VNPU3_3 port map (start_vn,clk,rst,Lc338,C218V338,C669V338,C1041V338,V338C218,V338C669,V338C1041,SI338,end_vn338);
V339:VNPU3_3 port map (start_vn,clk,rst,Lc339,C219V339,C670V339,C1042V339,V339C219,V339C670,V339C1042,SI339,end_vn339);
V340:VNPU3_3 port map (start_vn,clk,rst,Lc340,C220V340,C671V340,C1043V340,V340C220,V340C671,V340C1043,SI340,end_vn340);
V341:VNPU3_3 port map (start_vn,clk,rst,Lc341,C221V341,C672V341,C1044V341,V341C221,V341C672,V341C1044,SI341,end_vn341);
V342:VNPU3_3 port map (start_vn,clk,rst,Lc342,C222V342,C577V342,C1045V342,V342C222,V342C577,V342C1045,SI342,end_vn342);
V343:VNPU3_3 port map (start_vn,clk,rst,Lc343,C223V343,C578V343,C1046V343,V343C223,V343C578,V343C1046,SI343,end_vn343);
V344:VNPU3_3 port map (start_vn,clk,rst,Lc344,C224V344,C579V344,C1047V344,V344C224,V344C579,V344C1047,SI344,end_vn344);
V345:VNPU3_3 port map (start_vn,clk,rst,Lc345,C225V345,C580V345,C1048V345,V345C225,V345C580,V345C1048,SI345,end_vn345);
V346:VNPU3_3 port map (start_vn,clk,rst,Lc346,C226V346,C581V346,C1049V346,V346C226,V346C581,V346C1049,SI346,end_vn346);
V347:VNPU3_3 port map (start_vn,clk,rst,Lc347,C227V347,C582V347,C1050V347,V347C227,V347C582,V347C1050,SI347,end_vn347);
V348:VNPU3_3 port map (start_vn,clk,rst,Lc348,C228V348,C583V348,C1051V348,V348C228,V348C583,V348C1051,SI348,end_vn348);
V349:VNPU3_3 port map (start_vn,clk,rst,Lc349,C229V349,C584V349,C1052V349,V349C229,V349C584,V349C1052,SI349,end_vn349);
V350:VNPU3_3 port map (start_vn,clk,rst,Lc350,C230V350,C585V350,C1053V350,V350C230,V350C585,V350C1053,SI350,end_vn350);
V351:VNPU3_3 port map (start_vn,clk,rst,Lc351,C231V351,C586V351,C1054V351,V351C231,V351C586,V351C1054,SI351,end_vn351);
V352:VNPU3_3 port map (start_vn,clk,rst,Lc352,C232V352,C587V352,C1055V352,V352C232,V352C587,V352C1055,SI352,end_vn352);
V353:VNPU3_3 port map (start_vn,clk,rst,Lc353,C233V353,C588V353,C1056V353,V353C233,V353C588,V353C1056,SI353,end_vn353);
V354:VNPU3_3 port map (start_vn,clk,rst,Lc354,C234V354,C589V354,C961V354,V354C234,V354C589,V354C961,SI354,end_vn354);
V355:VNPU3_3 port map (start_vn,clk,rst,Lc355,C235V355,C590V355,C962V355,V355C235,V355C590,V355C962,SI355,end_vn355);
V356:VNPU3_3 port map (start_vn,clk,rst,Lc356,C236V356,C591V356,C963V356,V356C236,V356C591,V356C963,SI356,end_vn356);
V357:VNPU3_3 port map (start_vn,clk,rst,Lc357,C237V357,C592V357,C964V357,V357C237,V357C592,V357C964,SI357,end_vn357);
V358:VNPU3_3 port map (start_vn,clk,rst,Lc358,C238V358,C593V358,C965V358,V358C238,V358C593,V358C965,SI358,end_vn358);
V359:VNPU3_3 port map (start_vn,clk,rst,Lc359,C239V359,C594V359,C966V359,V359C239,V359C594,V359C966,SI359,end_vn359);
V360:VNPU3_3 port map (start_vn,clk,rst,Lc360,C240V360,C595V360,C967V360,V360C240,V360C595,V360C967,SI360,end_vn360);
V361:VNPU3_3 port map (start_vn,clk,rst,Lc361,C241V361,C596V361,C968V361,V361C241,V361C596,V361C968,SI361,end_vn361);
V362:VNPU3_3 port map (start_vn,clk,rst,Lc362,C242V362,C597V362,C969V362,V362C242,V362C597,V362C969,SI362,end_vn362);
V363:VNPU3_3 port map (start_vn,clk,rst,Lc363,C243V363,C598V363,C970V363,V363C243,V363C598,V363C970,SI363,end_vn363);
V364:VNPU3_3 port map (start_vn,clk,rst,Lc364,C244V364,C599V364,C971V364,V364C244,V364C599,V364C971,SI364,end_vn364);
V365:VNPU3_3 port map (start_vn,clk,rst,Lc365,C245V365,C600V365,C972V365,V365C245,V365C600,V365C972,SI365,end_vn365);
V366:VNPU3_3 port map (start_vn,clk,rst,Lc366,C246V366,C601V366,C973V366,V366C246,V366C601,V366C973,SI366,end_vn366);
V367:VNPU3_3 port map (start_vn,clk,rst,Lc367,C247V367,C602V367,C974V367,V367C247,V367C602,V367C974,SI367,end_vn367);
V368:VNPU3_3 port map (start_vn,clk,rst,Lc368,C248V368,C603V368,C975V368,V368C248,V368C603,V368C975,SI368,end_vn368);
V369:VNPU3_3 port map (start_vn,clk,rst,Lc369,C249V369,C604V369,C976V369,V369C249,V369C604,V369C976,SI369,end_vn369);
V370:VNPU3_3 port map (start_vn,clk,rst,Lc370,C250V370,C605V370,C977V370,V370C250,V370C605,V370C977,SI370,end_vn370);
V371:VNPU3_3 port map (start_vn,clk,rst,Lc371,C251V371,C606V371,C978V371,V371C251,V371C606,V371C978,SI371,end_vn371);
V372:VNPU3_3 port map (start_vn,clk,rst,Lc372,C252V372,C607V372,C979V372,V372C252,V372C607,V372C979,SI372,end_vn372);
V373:VNPU3_3 port map (start_vn,clk,rst,Lc373,C253V373,C608V373,C980V373,V373C253,V373C608,V373C980,SI373,end_vn373);
V374:VNPU3_3 port map (start_vn,clk,rst,Lc374,C254V374,C609V374,C981V374,V374C254,V374C609,V374C981,SI374,end_vn374);
V375:VNPU3_3 port map (start_vn,clk,rst,Lc375,C255V375,C610V375,C982V375,V375C255,V375C610,V375C982,SI375,end_vn375);
V376:VNPU3_3 port map (start_vn,clk,rst,Lc376,C256V376,C611V376,C983V376,V376C256,V376C611,V376C983,SI376,end_vn376);
V377:VNPU3_3 port map (start_vn,clk,rst,Lc377,C257V377,C612V377,C984V377,V377C257,V377C612,V377C984,SI377,end_vn377);
V378:VNPU3_3 port map (start_vn,clk,rst,Lc378,C258V378,C613V378,C985V378,V378C258,V378C613,V378C985,SI378,end_vn378);
V379:VNPU3_3 port map (start_vn,clk,rst,Lc379,C259V379,C614V379,C986V379,V379C259,V379C614,V379C986,SI379,end_vn379);
V380:VNPU3_3 port map (start_vn,clk,rst,Lc380,C260V380,C615V380,C987V380,V380C260,V380C615,V380C987,SI380,end_vn380);
V381:VNPU3_3 port map (start_vn,clk,rst,Lc381,C261V381,C616V381,C988V381,V381C261,V381C616,V381C988,SI381,end_vn381);
V382:VNPU3_3 port map (start_vn,clk,rst,Lc382,C262V382,C617V382,C989V382,V382C262,V382C617,V382C989,SI382,end_vn382);
V383:VNPU3_3 port map (start_vn,clk,rst,Lc383,C263V383,C618V383,C990V383,V383C263,V383C618,V383C990,SI383,end_vn383);
V384:VNPU3_3 port map (start_vn,clk,rst,Lc384,C264V384,C619V384,C991V384,V384C264,V384C619,V384C991,SI384,end_vn384);
V385:VNPU3_3 port map (start_vn,clk,rst,Lc385,C267V385,C531V385,C782V385,V385C267,V385C531,V385C782,SI385,end_vn385);
V386:VNPU3_3 port map (start_vn,clk,rst,Lc386,C268V386,C532V386,C783V386,V386C268,V386C532,V386C783,SI386,end_vn386);
V387:VNPU3_3 port map (start_vn,clk,rst,Lc387,C269V387,C533V387,C784V387,V387C269,V387C533,V387C784,SI387,end_vn387);
V388:VNPU3_3 port map (start_vn,clk,rst,Lc388,C270V388,C534V388,C785V388,V388C270,V388C534,V388C785,SI388,end_vn388);
V389:VNPU3_3 port map (start_vn,clk,rst,Lc389,C271V389,C535V389,C786V389,V389C271,V389C535,V389C786,SI389,end_vn389);
V390:VNPU3_3 port map (start_vn,clk,rst,Lc390,C272V390,C536V390,C787V390,V390C272,V390C536,V390C787,SI390,end_vn390);
V391:VNPU3_3 port map (start_vn,clk,rst,Lc391,C273V391,C537V391,C788V391,V391C273,V391C537,V391C788,SI391,end_vn391);
V392:VNPU3_3 port map (start_vn,clk,rst,Lc392,C274V392,C538V392,C789V392,V392C274,V392C538,V392C789,SI392,end_vn392);
V393:VNPU3_3 port map (start_vn,clk,rst,Lc393,C275V393,C539V393,C790V393,V393C275,V393C539,V393C790,SI393,end_vn393);
V394:VNPU3_3 port map (start_vn,clk,rst,Lc394,C276V394,C540V394,C791V394,V394C276,V394C540,V394C791,SI394,end_vn394);
V395:VNPU3_3 port map (start_vn,clk,rst,Lc395,C277V395,C541V395,C792V395,V395C277,V395C541,V395C792,SI395,end_vn395);
V396:VNPU3_3 port map (start_vn,clk,rst,Lc396,C278V396,C542V396,C793V396,V396C278,V396C542,V396C793,SI396,end_vn396);
V397:VNPU3_3 port map (start_vn,clk,rst,Lc397,C279V397,C543V397,C794V397,V397C279,V397C543,V397C794,SI397,end_vn397);
V398:VNPU3_3 port map (start_vn,clk,rst,Lc398,C280V398,C544V398,C795V398,V398C280,V398C544,V398C795,SI398,end_vn398);
V399:VNPU3_3 port map (start_vn,clk,rst,Lc399,C281V399,C545V399,C796V399,V399C281,V399C545,V399C796,SI399,end_vn399);
V400:VNPU3_3 port map (start_vn,clk,rst,Lc400,C282V400,C546V400,C797V400,V400C282,V400C546,V400C797,SI400,end_vn400);
V401:VNPU3_3 port map (start_vn,clk,rst,Lc401,C283V401,C547V401,C798V401,V401C283,V401C547,V401C798,SI401,end_vn401);
V402:VNPU3_3 port map (start_vn,clk,rst,Lc402,C284V402,C548V402,C799V402,V402C284,V402C548,V402C799,SI402,end_vn402);
V403:VNPU3_3 port map (start_vn,clk,rst,Lc403,C285V403,C549V403,C800V403,V403C285,V403C549,V403C800,SI403,end_vn403);
V404:VNPU3_3 port map (start_vn,clk,rst,Lc404,C286V404,C550V404,C801V404,V404C286,V404C550,V404C801,SI404,end_vn404);
V405:VNPU3_3 port map (start_vn,clk,rst,Lc405,C287V405,C551V405,C802V405,V405C287,V405C551,V405C802,SI405,end_vn405);
V406:VNPU3_3 port map (start_vn,clk,rst,Lc406,C288V406,C552V406,C803V406,V406C288,V406C552,V406C803,SI406,end_vn406);
V407:VNPU3_3 port map (start_vn,clk,rst,Lc407,C193V407,C553V407,C804V407,V407C193,V407C553,V407C804,SI407,end_vn407);
V408:VNPU3_3 port map (start_vn,clk,rst,Lc408,C194V408,C554V408,C805V408,V408C194,V408C554,V408C805,SI408,end_vn408);
V409:VNPU3_3 port map (start_vn,clk,rst,Lc409,C195V409,C555V409,C806V409,V409C195,V409C555,V409C806,SI409,end_vn409);
V410:VNPU3_3 port map (start_vn,clk,rst,Lc410,C196V410,C556V410,C807V410,V410C196,V410C556,V410C807,SI410,end_vn410);
V411:VNPU3_3 port map (start_vn,clk,rst,Lc411,C197V411,C557V411,C808V411,V411C197,V411C557,V411C808,SI411,end_vn411);
V412:VNPU3_3 port map (start_vn,clk,rst,Lc412,C198V412,C558V412,C809V412,V412C198,V412C558,V412C809,SI412,end_vn412);
V413:VNPU3_3 port map (start_vn,clk,rst,Lc413,C199V413,C559V413,C810V413,V413C199,V413C559,V413C810,SI413,end_vn413);
V414:VNPU3_3 port map (start_vn,clk,rst,Lc414,C200V414,C560V414,C811V414,V414C200,V414C560,V414C811,SI414,end_vn414);
V415:VNPU3_3 port map (start_vn,clk,rst,Lc415,C201V415,C561V415,C812V415,V415C201,V415C561,V415C812,SI415,end_vn415);
V416:VNPU3_3 port map (start_vn,clk,rst,Lc416,C202V416,C562V416,C813V416,V416C202,V416C562,V416C813,SI416,end_vn416);
V417:VNPU3_3 port map (start_vn,clk,rst,Lc417,C203V417,C563V417,C814V417,V417C203,V417C563,V417C814,SI417,end_vn417);
V418:VNPU3_3 port map (start_vn,clk,rst,Lc418,C204V418,C564V418,C815V418,V418C204,V418C564,V418C815,SI418,end_vn418);
V419:VNPU3_3 port map (start_vn,clk,rst,Lc419,C205V419,C565V419,C816V419,V419C205,V419C565,V419C816,SI419,end_vn419);
V420:VNPU3_3 port map (start_vn,clk,rst,Lc420,C206V420,C566V420,C817V420,V420C206,V420C566,V420C817,SI420,end_vn420);
V421:VNPU3_3 port map (start_vn,clk,rst,Lc421,C207V421,C567V421,C818V421,V421C207,V421C567,V421C818,SI421,end_vn421);
V422:VNPU3_3 port map (start_vn,clk,rst,Lc422,C208V422,C568V422,C819V422,V422C208,V422C568,V422C819,SI422,end_vn422);
V423:VNPU3_3 port map (start_vn,clk,rst,Lc423,C209V423,C569V423,C820V423,V423C209,V423C569,V423C820,SI423,end_vn423);
V424:VNPU3_3 port map (start_vn,clk,rst,Lc424,C210V424,C570V424,C821V424,V424C210,V424C570,V424C821,SI424,end_vn424);
V425:VNPU3_3 port map (start_vn,clk,rst,Lc425,C211V425,C571V425,C822V425,V425C211,V425C571,V425C822,SI425,end_vn425);
V426:VNPU3_3 port map (start_vn,clk,rst,Lc426,C212V426,C572V426,C823V426,V426C212,V426C572,V426C823,SI426,end_vn426);
V427:VNPU3_3 port map (start_vn,clk,rst,Lc427,C213V427,C573V427,C824V427,V427C213,V427C573,V427C824,SI427,end_vn427);
V428:VNPU3_3 port map (start_vn,clk,rst,Lc428,C214V428,C574V428,C825V428,V428C214,V428C574,V428C825,SI428,end_vn428);
V429:VNPU3_3 port map (start_vn,clk,rst,Lc429,C215V429,C575V429,C826V429,V429C215,V429C575,V429C826,SI429,end_vn429);
V430:VNPU3_3 port map (start_vn,clk,rst,Lc430,C216V430,C576V430,C827V430,V430C216,V430C576,V430C827,SI430,end_vn430);
V431:VNPU3_3 port map (start_vn,clk,rst,Lc431,C217V431,C481V431,C828V431,V431C217,V431C481,V431C828,SI431,end_vn431);
V432:VNPU3_3 port map (start_vn,clk,rst,Lc432,C218V432,C482V432,C829V432,V432C218,V432C482,V432C829,SI432,end_vn432);
V433:VNPU3_3 port map (start_vn,clk,rst,Lc433,C219V433,C483V433,C830V433,V433C219,V433C483,V433C830,SI433,end_vn433);
V434:VNPU3_3 port map (start_vn,clk,rst,Lc434,C220V434,C484V434,C831V434,V434C220,V434C484,V434C831,SI434,end_vn434);
V435:VNPU3_3 port map (start_vn,clk,rst,Lc435,C221V435,C485V435,C832V435,V435C221,V435C485,V435C832,SI435,end_vn435);
V436:VNPU3_3 port map (start_vn,clk,rst,Lc436,C222V436,C486V436,C833V436,V436C222,V436C486,V436C833,SI436,end_vn436);
V437:VNPU3_3 port map (start_vn,clk,rst,Lc437,C223V437,C487V437,C834V437,V437C223,V437C487,V437C834,SI437,end_vn437);
V438:VNPU3_3 port map (start_vn,clk,rst,Lc438,C224V438,C488V438,C835V438,V438C224,V438C488,V438C835,SI438,end_vn438);
V439:VNPU3_3 port map (start_vn,clk,rst,Lc439,C225V439,C489V439,C836V439,V439C225,V439C489,V439C836,SI439,end_vn439);
V440:VNPU3_3 port map (start_vn,clk,rst,Lc440,C226V440,C490V440,C837V440,V440C226,V440C490,V440C837,SI440,end_vn440);
V441:VNPU3_3 port map (start_vn,clk,rst,Lc441,C227V441,C491V441,C838V441,V441C227,V441C491,V441C838,SI441,end_vn441);
V442:VNPU3_3 port map (start_vn,clk,rst,Lc442,C228V442,C492V442,C839V442,V442C228,V442C492,V442C839,SI442,end_vn442);
V443:VNPU3_3 port map (start_vn,clk,rst,Lc443,C229V443,C493V443,C840V443,V443C229,V443C493,V443C840,SI443,end_vn443);
V444:VNPU3_3 port map (start_vn,clk,rst,Lc444,C230V444,C494V444,C841V444,V444C230,V444C494,V444C841,SI444,end_vn444);
V445:VNPU3_3 port map (start_vn,clk,rst,Lc445,C231V445,C495V445,C842V445,V445C231,V445C495,V445C842,SI445,end_vn445);
V446:VNPU3_3 port map (start_vn,clk,rst,Lc446,C232V446,C496V446,C843V446,V446C232,V446C496,V446C843,SI446,end_vn446);
V447:VNPU3_3 port map (start_vn,clk,rst,Lc447,C233V447,C497V447,C844V447,V447C233,V447C497,V447C844,SI447,end_vn447);
V448:VNPU3_3 port map (start_vn,clk,rst,Lc448,C234V448,C498V448,C845V448,V448C234,V448C498,V448C845,SI448,end_vn448);
V449:VNPU3_3 port map (start_vn,clk,rst,Lc449,C235V449,C499V449,C846V449,V449C235,V449C499,V449C846,SI449,end_vn449);
V450:VNPU3_3 port map (start_vn,clk,rst,Lc450,C236V450,C500V450,C847V450,V450C236,V450C500,V450C847,SI450,end_vn450);
V451:VNPU3_3 port map (start_vn,clk,rst,Lc451,C237V451,C501V451,C848V451,V451C237,V451C501,V451C848,SI451,end_vn451);
V452:VNPU3_3 port map (start_vn,clk,rst,Lc452,C238V452,C502V452,C849V452,V452C238,V452C502,V452C849,SI452,end_vn452);
V453:VNPU3_3 port map (start_vn,clk,rst,Lc453,C239V453,C503V453,C850V453,V453C239,V453C503,V453C850,SI453,end_vn453);
V454:VNPU3_3 port map (start_vn,clk,rst,Lc454,C240V454,C504V454,C851V454,V454C240,V454C504,V454C851,SI454,end_vn454);
V455:VNPU3_3 port map (start_vn,clk,rst,Lc455,C241V455,C505V455,C852V455,V455C241,V455C505,V455C852,SI455,end_vn455);
V456:VNPU3_3 port map (start_vn,clk,rst,Lc456,C242V456,C506V456,C853V456,V456C242,V456C506,V456C853,SI456,end_vn456);
V457:VNPU3_3 port map (start_vn,clk,rst,Lc457,C243V457,C507V457,C854V457,V457C243,V457C507,V457C854,SI457,end_vn457);
V458:VNPU3_3 port map (start_vn,clk,rst,Lc458,C244V458,C508V458,C855V458,V458C244,V458C508,V458C855,SI458,end_vn458);
V459:VNPU3_3 port map (start_vn,clk,rst,Lc459,C245V459,C509V459,C856V459,V459C245,V459C509,V459C856,SI459,end_vn459);
V460:VNPU3_3 port map (start_vn,clk,rst,Lc460,C246V460,C510V460,C857V460,V460C246,V460C510,V460C857,SI460,end_vn460);
V461:VNPU3_3 port map (start_vn,clk,rst,Lc461,C247V461,C511V461,C858V461,V461C247,V461C511,V461C858,SI461,end_vn461);
V462:VNPU3_3 port map (start_vn,clk,rst,Lc462,C248V462,C512V462,C859V462,V462C248,V462C512,V462C859,SI462,end_vn462);
V463:VNPU3_3 port map (start_vn,clk,rst,Lc463,C249V463,C513V463,C860V463,V463C249,V463C513,V463C860,SI463,end_vn463);
V464:VNPU3_3 port map (start_vn,clk,rst,Lc464,C250V464,C514V464,C861V464,V464C250,V464C514,V464C861,SI464,end_vn464);
V465:VNPU3_3 port map (start_vn,clk,rst,Lc465,C251V465,C515V465,C862V465,V465C251,V465C515,V465C862,SI465,end_vn465);
V466:VNPU3_3 port map (start_vn,clk,rst,Lc466,C252V466,C516V466,C863V466,V466C252,V466C516,V466C863,SI466,end_vn466);
V467:VNPU3_3 port map (start_vn,clk,rst,Lc467,C253V467,C517V467,C864V467,V467C253,V467C517,V467C864,SI467,end_vn467);
V468:VNPU3_3 port map (start_vn,clk,rst,Lc468,C254V468,C518V468,C769V468,V468C254,V468C518,V468C769,SI468,end_vn468);
V469:VNPU3_3 port map (start_vn,clk,rst,Lc469,C255V469,C519V469,C770V469,V469C255,V469C519,V469C770,SI469,end_vn469);
V470:VNPU3_3 port map (start_vn,clk,rst,Lc470,C256V470,C520V470,C771V470,V470C256,V470C520,V470C771,SI470,end_vn470);
V471:VNPU3_3 port map (start_vn,clk,rst,Lc471,C257V471,C521V471,C772V471,V471C257,V471C521,V471C772,SI471,end_vn471);
V472:VNPU3_3 port map (start_vn,clk,rst,Lc472,C258V472,C522V472,C773V472,V472C258,V472C522,V472C773,SI472,end_vn472);
V473:VNPU3_3 port map (start_vn,clk,rst,Lc473,C259V473,C523V473,C774V473,V473C259,V473C523,V473C774,SI473,end_vn473);
V474:VNPU3_3 port map (start_vn,clk,rst,Lc474,C260V474,C524V474,C775V474,V474C260,V474C524,V474C775,SI474,end_vn474);
V475:VNPU3_3 port map (start_vn,clk,rst,Lc475,C261V475,C525V475,C776V475,V475C261,V475C525,V475C776,SI475,end_vn475);
V476:VNPU3_3 port map (start_vn,clk,rst,Lc476,C262V476,C526V476,C777V476,V476C262,V476C526,V476C777,SI476,end_vn476);
V477:VNPU3_3 port map (start_vn,clk,rst,Lc477,C263V477,C527V477,C778V477,V477C263,V477C527,V477C778,SI477,end_vn477);
V478:VNPU3_3 port map (start_vn,clk,rst,Lc478,C264V478,C528V478,C779V478,V478C264,V478C528,V478C779,SI478,end_vn478);
V479:VNPU3_3 port map (start_vn,clk,rst,Lc479,C265V479,C529V479,C780V479,V479C265,V479C529,V479C780,SI479,end_vn479);
V480:VNPU3_3 port map (start_vn,clk,rst,Lc480,C266V480,C530V480,C781V480,V480C266,V480C530,V480C781,SI480,end_vn480);
V481:VNPU6_6 port map (start_vn,clk,rst,Lc481,C171V481,C208V481,C537V481,C841V481,C867V481,C1087V481,V481C171,V481C208,V481C537,V481C841,V481C867,V481C1087,SI481,end_vn481);
V482:VNPU6_6 port map (start_vn,clk,rst,Lc482,C172V482,C209V482,C538V482,C842V482,C868V482,C1088V482,V482C172,V482C209,V482C538,V482C842,V482C868,V482C1088,SI482,end_vn482);
V483:VNPU6_6 port map (start_vn,clk,rst,Lc483,C173V483,C210V483,C539V483,C843V483,C869V483,C1089V483,V483C173,V483C210,V483C539,V483C843,V483C869,V483C1089,SI483,end_vn483);
V484:VNPU6_6 port map (start_vn,clk,rst,Lc484,C174V484,C211V484,C540V484,C844V484,C870V484,C1090V484,V484C174,V484C211,V484C540,V484C844,V484C870,V484C1090,SI484,end_vn484);
V485:VNPU6_6 port map (start_vn,clk,rst,Lc485,C175V485,C212V485,C541V485,C845V485,C871V485,C1091V485,V485C175,V485C212,V485C541,V485C845,V485C871,V485C1091,SI485,end_vn485);
V486:VNPU6_6 port map (start_vn,clk,rst,Lc486,C176V486,C213V486,C542V486,C846V486,C872V486,C1092V486,V486C176,V486C213,V486C542,V486C846,V486C872,V486C1092,SI486,end_vn486);
V487:VNPU6_6 port map (start_vn,clk,rst,Lc487,C177V487,C214V487,C543V487,C847V487,C873V487,C1093V487,V487C177,V487C214,V487C543,V487C847,V487C873,V487C1093,SI487,end_vn487);
V488:VNPU6_6 port map (start_vn,clk,rst,Lc488,C178V488,C215V488,C544V488,C848V488,C874V488,C1094V488,V488C178,V488C215,V488C544,V488C848,V488C874,V488C1094,SI488,end_vn488);
V489:VNPU6_6 port map (start_vn,clk,rst,Lc489,C179V489,C216V489,C545V489,C849V489,C875V489,C1095V489,V489C179,V489C216,V489C545,V489C849,V489C875,V489C1095,SI489,end_vn489);
V490:VNPU6_6 port map (start_vn,clk,rst,Lc490,C180V490,C217V490,C546V490,C850V490,C876V490,C1096V490,V490C180,V490C217,V490C546,V490C850,V490C876,V490C1096,SI490,end_vn490);
V491:VNPU6_6 port map (start_vn,clk,rst,Lc491,C181V491,C218V491,C547V491,C851V491,C877V491,C1097V491,V491C181,V491C218,V491C547,V491C851,V491C877,V491C1097,SI491,end_vn491);
V492:VNPU6_6 port map (start_vn,clk,rst,Lc492,C182V492,C219V492,C548V492,C852V492,C878V492,C1098V492,V492C182,V492C219,V492C548,V492C852,V492C878,V492C1098,SI492,end_vn492);
V493:VNPU6_6 port map (start_vn,clk,rst,Lc493,C183V493,C220V493,C549V493,C853V493,C879V493,C1099V493,V493C183,V493C220,V493C549,V493C853,V493C879,V493C1099,SI493,end_vn493);
V494:VNPU6_6 port map (start_vn,clk,rst,Lc494,C184V494,C221V494,C550V494,C854V494,C880V494,C1100V494,V494C184,V494C221,V494C550,V494C854,V494C880,V494C1100,SI494,end_vn494);
V495:VNPU6_6 port map (start_vn,clk,rst,Lc495,C185V495,C222V495,C551V495,C855V495,C881V495,C1101V495,V495C185,V495C222,V495C551,V495C855,V495C881,V495C1101,SI495,end_vn495);
V496:VNPU6_6 port map (start_vn,clk,rst,Lc496,C186V496,C223V496,C552V496,C856V496,C882V496,C1102V496,V496C186,V496C223,V496C552,V496C856,V496C882,V496C1102,SI496,end_vn496);
V497:VNPU6_6 port map (start_vn,clk,rst,Lc497,C187V497,C224V497,C553V497,C857V497,C883V497,C1103V497,V497C187,V497C224,V497C553,V497C857,V497C883,V497C1103,SI497,end_vn497);
V498:VNPU6_6 port map (start_vn,clk,rst,Lc498,C188V498,C225V498,C554V498,C858V498,C884V498,C1104V498,V498C188,V498C225,V498C554,V498C858,V498C884,V498C1104,SI498,end_vn498);
V499:VNPU6_6 port map (start_vn,clk,rst,Lc499,C189V499,C226V499,C555V499,C859V499,C885V499,C1105V499,V499C189,V499C226,V499C555,V499C859,V499C885,V499C1105,SI499,end_vn499);
V500:VNPU6_6 port map (start_vn,clk,rst,Lc500,C190V500,C227V500,C556V500,C860V500,C886V500,C1106V500,V500C190,V500C227,V500C556,V500C860,V500C886,V500C1106,SI500,end_vn500);
V501:VNPU6_6 port map (start_vn,clk,rst,Lc501,C191V501,C228V501,C557V501,C861V501,C887V501,C1107V501,V501C191,V501C228,V501C557,V501C861,V501C887,V501C1107,SI501,end_vn501);
V502:VNPU6_6 port map (start_vn,clk,rst,Lc502,C192V502,C229V502,C558V502,C862V502,C888V502,C1108V502,V502C192,V502C229,V502C558,V502C862,V502C888,V502C1108,SI502,end_vn502);
V503:VNPU6_6 port map (start_vn,clk,rst,Lc503,C97V503,C230V503,C559V503,C863V503,C889V503,C1109V503,V503C97,V503C230,V503C559,V503C863,V503C889,V503C1109,SI503,end_vn503);
V504:VNPU6_6 port map (start_vn,clk,rst,Lc504,C98V504,C231V504,C560V504,C864V504,C890V504,C1110V504,V504C98,V504C231,V504C560,V504C864,V504C890,V504C1110,SI504,end_vn504);
V505:VNPU6_6 port map (start_vn,clk,rst,Lc505,C99V505,C232V505,C561V505,C769V505,C891V505,C1111V505,V505C99,V505C232,V505C561,V505C769,V505C891,V505C1111,SI505,end_vn505);
V506:VNPU6_6 port map (start_vn,clk,rst,Lc506,C100V506,C233V506,C562V506,C770V506,C892V506,C1112V506,V506C100,V506C233,V506C562,V506C770,V506C892,V506C1112,SI506,end_vn506);
V507:VNPU6_6 port map (start_vn,clk,rst,Lc507,C101V507,C234V507,C563V507,C771V507,C893V507,C1113V507,V507C101,V507C234,V507C563,V507C771,V507C893,V507C1113,SI507,end_vn507);
V508:VNPU6_6 port map (start_vn,clk,rst,Lc508,C102V508,C235V508,C564V508,C772V508,C894V508,C1114V508,V508C102,V508C235,V508C564,V508C772,V508C894,V508C1114,SI508,end_vn508);
V509:VNPU6_6 port map (start_vn,clk,rst,Lc509,C103V509,C236V509,C565V509,C773V509,C895V509,C1115V509,V509C103,V509C236,V509C565,V509C773,V509C895,V509C1115,SI509,end_vn509);
V510:VNPU6_6 port map (start_vn,clk,rst,Lc510,C104V510,C237V510,C566V510,C774V510,C896V510,C1116V510,V510C104,V510C237,V510C566,V510C774,V510C896,V510C1116,SI510,end_vn510);
V511:VNPU6_6 port map (start_vn,clk,rst,Lc511,C105V511,C238V511,C567V511,C775V511,C897V511,C1117V511,V511C105,V511C238,V511C567,V511C775,V511C897,V511C1117,SI511,end_vn511);
V512:VNPU6_6 port map (start_vn,clk,rst,Lc512,C106V512,C239V512,C568V512,C776V512,C898V512,C1118V512,V512C106,V512C239,V512C568,V512C776,V512C898,V512C1118,SI512,end_vn512);
V513:VNPU6_6 port map (start_vn,clk,rst,Lc513,C107V513,C240V513,C569V513,C777V513,C899V513,C1119V513,V513C107,V513C240,V513C569,V513C777,V513C899,V513C1119,SI513,end_vn513);
V514:VNPU6_6 port map (start_vn,clk,rst,Lc514,C108V514,C241V514,C570V514,C778V514,C900V514,C1120V514,V514C108,V514C241,V514C570,V514C778,V514C900,V514C1120,SI514,end_vn514);
V515:VNPU6_6 port map (start_vn,clk,rst,Lc515,C109V515,C242V515,C571V515,C779V515,C901V515,C1121V515,V515C109,V515C242,V515C571,V515C779,V515C901,V515C1121,SI515,end_vn515);
V516:VNPU6_6 port map (start_vn,clk,rst,Lc516,C110V516,C243V516,C572V516,C780V516,C902V516,C1122V516,V516C110,V516C243,V516C572,V516C780,V516C902,V516C1122,SI516,end_vn516);
V517:VNPU6_6 port map (start_vn,clk,rst,Lc517,C111V517,C244V517,C573V517,C781V517,C903V517,C1123V517,V517C111,V517C244,V517C573,V517C781,V517C903,V517C1123,SI517,end_vn517);
V518:VNPU6_6 port map (start_vn,clk,rst,Lc518,C112V518,C245V518,C574V518,C782V518,C904V518,C1124V518,V518C112,V518C245,V518C574,V518C782,V518C904,V518C1124,SI518,end_vn518);
V519:VNPU6_6 port map (start_vn,clk,rst,Lc519,C113V519,C246V519,C575V519,C783V519,C905V519,C1125V519,V519C113,V519C246,V519C575,V519C783,V519C905,V519C1125,SI519,end_vn519);
V520:VNPU6_6 port map (start_vn,clk,rst,Lc520,C114V520,C247V520,C576V520,C784V520,C906V520,C1126V520,V520C114,V520C247,V520C576,V520C784,V520C906,V520C1126,SI520,end_vn520);
V521:VNPU6_6 port map (start_vn,clk,rst,Lc521,C115V521,C248V521,C481V521,C785V521,C907V521,C1127V521,V521C115,V521C248,V521C481,V521C785,V521C907,V521C1127,SI521,end_vn521);
V522:VNPU6_6 port map (start_vn,clk,rst,Lc522,C116V522,C249V522,C482V522,C786V522,C908V522,C1128V522,V522C116,V522C249,V522C482,V522C786,V522C908,V522C1128,SI522,end_vn522);
V523:VNPU6_6 port map (start_vn,clk,rst,Lc523,C117V523,C250V523,C483V523,C787V523,C909V523,C1129V523,V523C117,V523C250,V523C483,V523C787,V523C909,V523C1129,SI523,end_vn523);
V524:VNPU6_6 port map (start_vn,clk,rst,Lc524,C118V524,C251V524,C484V524,C788V524,C910V524,C1130V524,V524C118,V524C251,V524C484,V524C788,V524C910,V524C1130,SI524,end_vn524);
V525:VNPU6_6 port map (start_vn,clk,rst,Lc525,C119V525,C252V525,C485V525,C789V525,C911V525,C1131V525,V525C119,V525C252,V525C485,V525C789,V525C911,V525C1131,SI525,end_vn525);
V526:VNPU6_6 port map (start_vn,clk,rst,Lc526,C120V526,C253V526,C486V526,C790V526,C912V526,C1132V526,V526C120,V526C253,V526C486,V526C790,V526C912,V526C1132,SI526,end_vn526);
V527:VNPU6_6 port map (start_vn,clk,rst,Lc527,C121V527,C254V527,C487V527,C791V527,C913V527,C1133V527,V527C121,V527C254,V527C487,V527C791,V527C913,V527C1133,SI527,end_vn527);
V528:VNPU6_6 port map (start_vn,clk,rst,Lc528,C122V528,C255V528,C488V528,C792V528,C914V528,C1134V528,V528C122,V528C255,V528C488,V528C792,V528C914,V528C1134,SI528,end_vn528);
V529:VNPU6_6 port map (start_vn,clk,rst,Lc529,C123V529,C256V529,C489V529,C793V529,C915V529,C1135V529,V529C123,V529C256,V529C489,V529C793,V529C915,V529C1135,SI529,end_vn529);
V530:VNPU6_6 port map (start_vn,clk,rst,Lc530,C124V530,C257V530,C490V530,C794V530,C916V530,C1136V530,V530C124,V530C257,V530C490,V530C794,V530C916,V530C1136,SI530,end_vn530);
V531:VNPU6_6 port map (start_vn,clk,rst,Lc531,C125V531,C258V531,C491V531,C795V531,C917V531,C1137V531,V531C125,V531C258,V531C491,V531C795,V531C917,V531C1137,SI531,end_vn531);
V532:VNPU6_6 port map (start_vn,clk,rst,Lc532,C126V532,C259V532,C492V532,C796V532,C918V532,C1138V532,V532C126,V532C259,V532C492,V532C796,V532C918,V532C1138,SI532,end_vn532);
V533:VNPU6_6 port map (start_vn,clk,rst,Lc533,C127V533,C260V533,C493V533,C797V533,C919V533,C1139V533,V533C127,V533C260,V533C493,V533C797,V533C919,V533C1139,SI533,end_vn533);
V534:VNPU6_6 port map (start_vn,clk,rst,Lc534,C128V534,C261V534,C494V534,C798V534,C920V534,C1140V534,V534C128,V534C261,V534C494,V534C798,V534C920,V534C1140,SI534,end_vn534);
V535:VNPU6_6 port map (start_vn,clk,rst,Lc535,C129V535,C262V535,C495V535,C799V535,C921V535,C1141V535,V535C129,V535C262,V535C495,V535C799,V535C921,V535C1141,SI535,end_vn535);
V536:VNPU6_6 port map (start_vn,clk,rst,Lc536,C130V536,C263V536,C496V536,C800V536,C922V536,C1142V536,V536C130,V536C263,V536C496,V536C800,V536C922,V536C1142,SI536,end_vn536);
V537:VNPU6_6 port map (start_vn,clk,rst,Lc537,C131V537,C264V537,C497V537,C801V537,C923V537,C1143V537,V537C131,V537C264,V537C497,V537C801,V537C923,V537C1143,SI537,end_vn537);
V538:VNPU6_6 port map (start_vn,clk,rst,Lc538,C132V538,C265V538,C498V538,C802V538,C924V538,C1144V538,V538C132,V538C265,V538C498,V538C802,V538C924,V538C1144,SI538,end_vn538);
V539:VNPU6_6 port map (start_vn,clk,rst,Lc539,C133V539,C266V539,C499V539,C803V539,C925V539,C1145V539,V539C133,V539C266,V539C499,V539C803,V539C925,V539C1145,SI539,end_vn539);
V540:VNPU6_6 port map (start_vn,clk,rst,Lc540,C134V540,C267V540,C500V540,C804V540,C926V540,C1146V540,V540C134,V540C267,V540C500,V540C804,V540C926,V540C1146,SI540,end_vn540);
V541:VNPU6_6 port map (start_vn,clk,rst,Lc541,C135V541,C268V541,C501V541,C805V541,C927V541,C1147V541,V541C135,V541C268,V541C501,V541C805,V541C927,V541C1147,SI541,end_vn541);
V542:VNPU6_6 port map (start_vn,clk,rst,Lc542,C136V542,C269V542,C502V542,C806V542,C928V542,C1148V542,V542C136,V542C269,V542C502,V542C806,V542C928,V542C1148,SI542,end_vn542);
V543:VNPU6_6 port map (start_vn,clk,rst,Lc543,C137V543,C270V543,C503V543,C807V543,C929V543,C1149V543,V543C137,V543C270,V543C503,V543C807,V543C929,V543C1149,SI543,end_vn543);
V544:VNPU6_6 port map (start_vn,clk,rst,Lc544,C138V544,C271V544,C504V544,C808V544,C930V544,C1150V544,V544C138,V544C271,V544C504,V544C808,V544C930,V544C1150,SI544,end_vn544);
V545:VNPU6_6 port map (start_vn,clk,rst,Lc545,C139V545,C272V545,C505V545,C809V545,C931V545,C1151V545,V545C139,V545C272,V545C505,V545C809,V545C931,V545C1151,SI545,end_vn545);
V546:VNPU6_6 port map (start_vn,clk,rst,Lc546,C140V546,C273V546,C506V546,C810V546,C932V546,C1152V546,V546C140,V546C273,V546C506,V546C810,V546C932,V546C1152,SI546,end_vn546);
V547:VNPU6_6 port map (start_vn,clk,rst,Lc547,C141V547,C274V547,C507V547,C811V547,C933V547,C1057V547,V547C141,V547C274,V547C507,V547C811,V547C933,V547C1057,SI547,end_vn547);
V548:VNPU6_6 port map (start_vn,clk,rst,Lc548,C142V548,C275V548,C508V548,C812V548,C934V548,C1058V548,V548C142,V548C275,V548C508,V548C812,V548C934,V548C1058,SI548,end_vn548);
V549:VNPU6_6 port map (start_vn,clk,rst,Lc549,C143V549,C276V549,C509V549,C813V549,C935V549,C1059V549,V549C143,V549C276,V549C509,V549C813,V549C935,V549C1059,SI549,end_vn549);
V550:VNPU6_6 port map (start_vn,clk,rst,Lc550,C144V550,C277V550,C510V550,C814V550,C936V550,C1060V550,V550C144,V550C277,V550C510,V550C814,V550C936,V550C1060,SI550,end_vn550);
V551:VNPU6_6 port map (start_vn,clk,rst,Lc551,C145V551,C278V551,C511V551,C815V551,C937V551,C1061V551,V551C145,V551C278,V551C511,V551C815,V551C937,V551C1061,SI551,end_vn551);
V552:VNPU6_6 port map (start_vn,clk,rst,Lc552,C146V552,C279V552,C512V552,C816V552,C938V552,C1062V552,V552C146,V552C279,V552C512,V552C816,V552C938,V552C1062,SI552,end_vn552);
V553:VNPU6_6 port map (start_vn,clk,rst,Lc553,C147V553,C280V553,C513V553,C817V553,C939V553,C1063V553,V553C147,V553C280,V553C513,V553C817,V553C939,V553C1063,SI553,end_vn553);
V554:VNPU6_6 port map (start_vn,clk,rst,Lc554,C148V554,C281V554,C514V554,C818V554,C940V554,C1064V554,V554C148,V554C281,V554C514,V554C818,V554C940,V554C1064,SI554,end_vn554);
V555:VNPU6_6 port map (start_vn,clk,rst,Lc555,C149V555,C282V555,C515V555,C819V555,C941V555,C1065V555,V555C149,V555C282,V555C515,V555C819,V555C941,V555C1065,SI555,end_vn555);
V556:VNPU6_6 port map (start_vn,clk,rst,Lc556,C150V556,C283V556,C516V556,C820V556,C942V556,C1066V556,V556C150,V556C283,V556C516,V556C820,V556C942,V556C1066,SI556,end_vn556);
V557:VNPU6_6 port map (start_vn,clk,rst,Lc557,C151V557,C284V557,C517V557,C821V557,C943V557,C1067V557,V557C151,V557C284,V557C517,V557C821,V557C943,V557C1067,SI557,end_vn557);
V558:VNPU6_6 port map (start_vn,clk,rst,Lc558,C152V558,C285V558,C518V558,C822V558,C944V558,C1068V558,V558C152,V558C285,V558C518,V558C822,V558C944,V558C1068,SI558,end_vn558);
V559:VNPU6_6 port map (start_vn,clk,rst,Lc559,C153V559,C286V559,C519V559,C823V559,C945V559,C1069V559,V559C153,V559C286,V559C519,V559C823,V559C945,V559C1069,SI559,end_vn559);
V560:VNPU6_6 port map (start_vn,clk,rst,Lc560,C154V560,C287V560,C520V560,C824V560,C946V560,C1070V560,V560C154,V560C287,V560C520,V560C824,V560C946,V560C1070,SI560,end_vn560);
V561:VNPU6_6 port map (start_vn,clk,rst,Lc561,C155V561,C288V561,C521V561,C825V561,C947V561,C1071V561,V561C155,V561C288,V561C521,V561C825,V561C947,V561C1071,SI561,end_vn561);
V562:VNPU6_6 port map (start_vn,clk,rst,Lc562,C156V562,C193V562,C522V562,C826V562,C948V562,C1072V562,V562C156,V562C193,V562C522,V562C826,V562C948,V562C1072,SI562,end_vn562);
V563:VNPU6_6 port map (start_vn,clk,rst,Lc563,C157V563,C194V563,C523V563,C827V563,C949V563,C1073V563,V563C157,V563C194,V563C523,V563C827,V563C949,V563C1073,SI563,end_vn563);
V564:VNPU6_6 port map (start_vn,clk,rst,Lc564,C158V564,C195V564,C524V564,C828V564,C950V564,C1074V564,V564C158,V564C195,V564C524,V564C828,V564C950,V564C1074,SI564,end_vn564);
V565:VNPU6_6 port map (start_vn,clk,rst,Lc565,C159V565,C196V565,C525V565,C829V565,C951V565,C1075V565,V565C159,V565C196,V565C525,V565C829,V565C951,V565C1075,SI565,end_vn565);
V566:VNPU6_6 port map (start_vn,clk,rst,Lc566,C160V566,C197V566,C526V566,C830V566,C952V566,C1076V566,V566C160,V566C197,V566C526,V566C830,V566C952,V566C1076,SI566,end_vn566);
V567:VNPU6_6 port map (start_vn,clk,rst,Lc567,C161V567,C198V567,C527V567,C831V567,C953V567,C1077V567,V567C161,V567C198,V567C527,V567C831,V567C953,V567C1077,SI567,end_vn567);
V568:VNPU6_6 port map (start_vn,clk,rst,Lc568,C162V568,C199V568,C528V568,C832V568,C954V568,C1078V568,V568C162,V568C199,V568C528,V568C832,V568C954,V568C1078,SI568,end_vn568);
V569:VNPU6_6 port map (start_vn,clk,rst,Lc569,C163V569,C200V569,C529V569,C833V569,C955V569,C1079V569,V569C163,V569C200,V569C529,V569C833,V569C955,V569C1079,SI569,end_vn569);
V570:VNPU6_6 port map (start_vn,clk,rst,Lc570,C164V570,C201V570,C530V570,C834V570,C956V570,C1080V570,V570C164,V570C201,V570C530,V570C834,V570C956,V570C1080,SI570,end_vn570);
V571:VNPU6_6 port map (start_vn,clk,rst,Lc571,C165V571,C202V571,C531V571,C835V571,C957V571,C1081V571,V571C165,V571C202,V571C531,V571C835,V571C957,V571C1081,SI571,end_vn571);
V572:VNPU6_6 port map (start_vn,clk,rst,Lc572,C166V572,C203V572,C532V572,C836V572,C958V572,C1082V572,V572C166,V572C203,V572C532,V572C836,V572C958,V572C1082,SI572,end_vn572);
V573:VNPU6_6 port map (start_vn,clk,rst,Lc573,C167V573,C204V573,C533V573,C837V573,C959V573,C1083V573,V573C167,V573C204,V573C533,V573C837,V573C959,V573C1083,SI573,end_vn573);
V574:VNPU6_6 port map (start_vn,clk,rst,Lc574,C168V574,C205V574,C534V574,C838V574,C960V574,C1084V574,V574C168,V574C205,V574C534,V574C838,V574C960,V574C1084,SI574,end_vn574);
V575:VNPU6_6 port map (start_vn,clk,rst,Lc575,C169V575,C206V575,C535V575,C839V575,C865V575,C1085V575,V575C169,V575C206,V575C535,V575C839,V575C865,V575C1085,SI575,end_vn575);
V576:VNPU6_6 port map (start_vn,clk,rst,Lc576,C170V576,C207V576,C536V576,C840V576,C866V576,C1086V576,V576C170,V576C207,V576C536,V576C840,V576C866,V576C1086,SI576,end_vn576);
V577:VNPU3_3 port map (start_vn,clk,rst,Lc577,C114V577,C397V577,C767V577,V577C114,V577C397,V577C767,SI577,end_vn577);
V578:VNPU3_3 port map (start_vn,clk,rst,Lc578,C115V578,C398V578,C768V578,V578C115,V578C398,V578C768,SI578,end_vn578);
V579:VNPU3_3 port map (start_vn,clk,rst,Lc579,C116V579,C399V579,C673V579,V579C116,V579C399,V579C673,SI579,end_vn579);
V580:VNPU3_3 port map (start_vn,clk,rst,Lc580,C117V580,C400V580,C674V580,V580C117,V580C400,V580C674,SI580,end_vn580);
V581:VNPU3_3 port map (start_vn,clk,rst,Lc581,C118V581,C401V581,C675V581,V581C118,V581C401,V581C675,SI581,end_vn581);
V582:VNPU3_3 port map (start_vn,clk,rst,Lc582,C119V582,C402V582,C676V582,V582C119,V582C402,V582C676,SI582,end_vn582);
V583:VNPU3_3 port map (start_vn,clk,rst,Lc583,C120V583,C403V583,C677V583,V583C120,V583C403,V583C677,SI583,end_vn583);
V584:VNPU3_3 port map (start_vn,clk,rst,Lc584,C121V584,C404V584,C678V584,V584C121,V584C404,V584C678,SI584,end_vn584);
V585:VNPU3_3 port map (start_vn,clk,rst,Lc585,C122V585,C405V585,C679V585,V585C122,V585C405,V585C679,SI585,end_vn585);
V586:VNPU3_3 port map (start_vn,clk,rst,Lc586,C123V586,C406V586,C680V586,V586C123,V586C406,V586C680,SI586,end_vn586);
V587:VNPU3_3 port map (start_vn,clk,rst,Lc587,C124V587,C407V587,C681V587,V587C124,V587C407,V587C681,SI587,end_vn587);
V588:VNPU3_3 port map (start_vn,clk,rst,Lc588,C125V588,C408V588,C682V588,V588C125,V588C408,V588C682,SI588,end_vn588);
V589:VNPU3_3 port map (start_vn,clk,rst,Lc589,C126V589,C409V589,C683V589,V589C126,V589C409,V589C683,SI589,end_vn589);
V590:VNPU3_3 port map (start_vn,clk,rst,Lc590,C127V590,C410V590,C684V590,V590C127,V590C410,V590C684,SI590,end_vn590);
V591:VNPU3_3 port map (start_vn,clk,rst,Lc591,C128V591,C411V591,C685V591,V591C128,V591C411,V591C685,SI591,end_vn591);
V592:VNPU3_3 port map (start_vn,clk,rst,Lc592,C129V592,C412V592,C686V592,V592C129,V592C412,V592C686,SI592,end_vn592);
V593:VNPU3_3 port map (start_vn,clk,rst,Lc593,C130V593,C413V593,C687V593,V593C130,V593C413,V593C687,SI593,end_vn593);
V594:VNPU3_3 port map (start_vn,clk,rst,Lc594,C131V594,C414V594,C688V594,V594C131,V594C414,V594C688,SI594,end_vn594);
V595:VNPU3_3 port map (start_vn,clk,rst,Lc595,C132V595,C415V595,C689V595,V595C132,V595C415,V595C689,SI595,end_vn595);
V596:VNPU3_3 port map (start_vn,clk,rst,Lc596,C133V596,C416V596,C690V596,V596C133,V596C416,V596C690,SI596,end_vn596);
V597:VNPU3_3 port map (start_vn,clk,rst,Lc597,C134V597,C417V597,C691V597,V597C134,V597C417,V597C691,SI597,end_vn597);
V598:VNPU3_3 port map (start_vn,clk,rst,Lc598,C135V598,C418V598,C692V598,V598C135,V598C418,V598C692,SI598,end_vn598);
V599:VNPU3_3 port map (start_vn,clk,rst,Lc599,C136V599,C419V599,C693V599,V599C136,V599C419,V599C693,SI599,end_vn599);
V600:VNPU3_3 port map (start_vn,clk,rst,Lc600,C137V600,C420V600,C694V600,V600C137,V600C420,V600C694,SI600,end_vn600);
V601:VNPU3_3 port map (start_vn,clk,rst,Lc601,C138V601,C421V601,C695V601,V601C138,V601C421,V601C695,SI601,end_vn601);
V602:VNPU3_3 port map (start_vn,clk,rst,Lc602,C139V602,C422V602,C696V602,V602C139,V602C422,V602C696,SI602,end_vn602);
V603:VNPU3_3 port map (start_vn,clk,rst,Lc603,C140V603,C423V603,C697V603,V603C140,V603C423,V603C697,SI603,end_vn603);
V604:VNPU3_3 port map (start_vn,clk,rst,Lc604,C141V604,C424V604,C698V604,V604C141,V604C424,V604C698,SI604,end_vn604);
V605:VNPU3_3 port map (start_vn,clk,rst,Lc605,C142V605,C425V605,C699V605,V605C142,V605C425,V605C699,SI605,end_vn605);
V606:VNPU3_3 port map (start_vn,clk,rst,Lc606,C143V606,C426V606,C700V606,V606C143,V606C426,V606C700,SI606,end_vn606);
V607:VNPU3_3 port map (start_vn,clk,rst,Lc607,C144V607,C427V607,C701V607,V607C144,V607C427,V607C701,SI607,end_vn607);
V608:VNPU3_3 port map (start_vn,clk,rst,Lc608,C145V608,C428V608,C702V608,V608C145,V608C428,V608C702,SI608,end_vn608);
V609:VNPU3_3 port map (start_vn,clk,rst,Lc609,C146V609,C429V609,C703V609,V609C146,V609C429,V609C703,SI609,end_vn609);
V610:VNPU3_3 port map (start_vn,clk,rst,Lc610,C147V610,C430V610,C704V610,V610C147,V610C430,V610C704,SI610,end_vn610);
V611:VNPU3_3 port map (start_vn,clk,rst,Lc611,C148V611,C431V611,C705V611,V611C148,V611C431,V611C705,SI611,end_vn611);
V612:VNPU3_3 port map (start_vn,clk,rst,Lc612,C149V612,C432V612,C706V612,V612C149,V612C432,V612C706,SI612,end_vn612);
V613:VNPU3_3 port map (start_vn,clk,rst,Lc613,C150V613,C433V613,C707V613,V613C150,V613C433,V613C707,SI613,end_vn613);
V614:VNPU3_3 port map (start_vn,clk,rst,Lc614,C151V614,C434V614,C708V614,V614C151,V614C434,V614C708,SI614,end_vn614);
V615:VNPU3_3 port map (start_vn,clk,rst,Lc615,C152V615,C435V615,C709V615,V615C152,V615C435,V615C709,SI615,end_vn615);
V616:VNPU3_3 port map (start_vn,clk,rst,Lc616,C153V616,C436V616,C710V616,V616C153,V616C436,V616C710,SI616,end_vn616);
V617:VNPU3_3 port map (start_vn,clk,rst,Lc617,C154V617,C437V617,C711V617,V617C154,V617C437,V617C711,SI617,end_vn617);
V618:VNPU3_3 port map (start_vn,clk,rst,Lc618,C155V618,C438V618,C712V618,V618C155,V618C438,V618C712,SI618,end_vn618);
V619:VNPU3_3 port map (start_vn,clk,rst,Lc619,C156V619,C439V619,C713V619,V619C156,V619C439,V619C713,SI619,end_vn619);
V620:VNPU3_3 port map (start_vn,clk,rst,Lc620,C157V620,C440V620,C714V620,V620C157,V620C440,V620C714,SI620,end_vn620);
V621:VNPU3_3 port map (start_vn,clk,rst,Lc621,C158V621,C441V621,C715V621,V621C158,V621C441,V621C715,SI621,end_vn621);
V622:VNPU3_3 port map (start_vn,clk,rst,Lc622,C159V622,C442V622,C716V622,V622C159,V622C442,V622C716,SI622,end_vn622);
V623:VNPU3_3 port map (start_vn,clk,rst,Lc623,C160V623,C443V623,C717V623,V623C160,V623C443,V623C717,SI623,end_vn623);
V624:VNPU3_3 port map (start_vn,clk,rst,Lc624,C161V624,C444V624,C718V624,V624C161,V624C444,V624C718,SI624,end_vn624);
V625:VNPU3_3 port map (start_vn,clk,rst,Lc625,C162V625,C445V625,C719V625,V625C162,V625C445,V625C719,SI625,end_vn625);
V626:VNPU3_3 port map (start_vn,clk,rst,Lc626,C163V626,C446V626,C720V626,V626C163,V626C446,V626C720,SI626,end_vn626);
V627:VNPU3_3 port map (start_vn,clk,rst,Lc627,C164V627,C447V627,C721V627,V627C164,V627C447,V627C721,SI627,end_vn627);
V628:VNPU3_3 port map (start_vn,clk,rst,Lc628,C165V628,C448V628,C722V628,V628C165,V628C448,V628C722,SI628,end_vn628);
V629:VNPU3_3 port map (start_vn,clk,rst,Lc629,C166V629,C449V629,C723V629,V629C166,V629C449,V629C723,SI629,end_vn629);
V630:VNPU3_3 port map (start_vn,clk,rst,Lc630,C167V630,C450V630,C724V630,V630C167,V630C450,V630C724,SI630,end_vn630);
V631:VNPU3_3 port map (start_vn,clk,rst,Lc631,C168V631,C451V631,C725V631,V631C168,V631C451,V631C725,SI631,end_vn631);
V632:VNPU3_3 port map (start_vn,clk,rst,Lc632,C169V632,C452V632,C726V632,V632C169,V632C452,V632C726,SI632,end_vn632);
V633:VNPU3_3 port map (start_vn,clk,rst,Lc633,C170V633,C453V633,C727V633,V633C170,V633C453,V633C727,SI633,end_vn633);
V634:VNPU3_3 port map (start_vn,clk,rst,Lc634,C171V634,C454V634,C728V634,V634C171,V634C454,V634C728,SI634,end_vn634);
V635:VNPU3_3 port map (start_vn,clk,rst,Lc635,C172V635,C455V635,C729V635,V635C172,V635C455,V635C729,SI635,end_vn635);
V636:VNPU3_3 port map (start_vn,clk,rst,Lc636,C173V636,C456V636,C730V636,V636C173,V636C456,V636C730,SI636,end_vn636);
V637:VNPU3_3 port map (start_vn,clk,rst,Lc637,C174V637,C457V637,C731V637,V637C174,V637C457,V637C731,SI637,end_vn637);
V638:VNPU3_3 port map (start_vn,clk,rst,Lc638,C175V638,C458V638,C732V638,V638C175,V638C458,V638C732,SI638,end_vn638);
V639:VNPU3_3 port map (start_vn,clk,rst,Lc639,C176V639,C459V639,C733V639,V639C176,V639C459,V639C733,SI639,end_vn639);
V640:VNPU3_3 port map (start_vn,clk,rst,Lc640,C177V640,C460V640,C734V640,V640C177,V640C460,V640C734,SI640,end_vn640);
V641:VNPU3_3 port map (start_vn,clk,rst,Lc641,C178V641,C461V641,C735V641,V641C178,V641C461,V641C735,SI641,end_vn641);
V642:VNPU3_3 port map (start_vn,clk,rst,Lc642,C179V642,C462V642,C736V642,V642C179,V642C462,V642C736,SI642,end_vn642);
V643:VNPU3_3 port map (start_vn,clk,rst,Lc643,C180V643,C463V643,C737V643,V643C180,V643C463,V643C737,SI643,end_vn643);
V644:VNPU3_3 port map (start_vn,clk,rst,Lc644,C181V644,C464V644,C738V644,V644C181,V644C464,V644C738,SI644,end_vn644);
V645:VNPU3_3 port map (start_vn,clk,rst,Lc645,C182V645,C465V645,C739V645,V645C182,V645C465,V645C739,SI645,end_vn645);
V646:VNPU3_3 port map (start_vn,clk,rst,Lc646,C183V646,C466V646,C740V646,V646C183,V646C466,V646C740,SI646,end_vn646);
V647:VNPU3_3 port map (start_vn,clk,rst,Lc647,C184V647,C467V647,C741V647,V647C184,V647C467,V647C741,SI647,end_vn647);
V648:VNPU3_3 port map (start_vn,clk,rst,Lc648,C185V648,C468V648,C742V648,V648C185,V648C468,V648C742,SI648,end_vn648);
V649:VNPU3_3 port map (start_vn,clk,rst,Lc649,C186V649,C469V649,C743V649,V649C186,V649C469,V649C743,SI649,end_vn649);
V650:VNPU3_3 port map (start_vn,clk,rst,Lc650,C187V650,C470V650,C744V650,V650C187,V650C470,V650C744,SI650,end_vn650);
V651:VNPU3_3 port map (start_vn,clk,rst,Lc651,C188V651,C471V651,C745V651,V651C188,V651C471,V651C745,SI651,end_vn651);
V652:VNPU3_3 port map (start_vn,clk,rst,Lc652,C189V652,C472V652,C746V652,V652C189,V652C472,V652C746,SI652,end_vn652);
V653:VNPU3_3 port map (start_vn,clk,rst,Lc653,C190V653,C473V653,C747V653,V653C190,V653C473,V653C747,SI653,end_vn653);
V654:VNPU3_3 port map (start_vn,clk,rst,Lc654,C191V654,C474V654,C748V654,V654C191,V654C474,V654C748,SI654,end_vn654);
V655:VNPU3_3 port map (start_vn,clk,rst,Lc655,C192V655,C475V655,C749V655,V655C192,V655C475,V655C749,SI655,end_vn655);
V656:VNPU3_3 port map (start_vn,clk,rst,Lc656,C97V656,C476V656,C750V656,V656C97,V656C476,V656C750,SI656,end_vn656);
V657:VNPU3_3 port map (start_vn,clk,rst,Lc657,C98V657,C477V657,C751V657,V657C98,V657C477,V657C751,SI657,end_vn657);
V658:VNPU3_3 port map (start_vn,clk,rst,Lc658,C99V658,C478V658,C752V658,V658C99,V658C478,V658C752,SI658,end_vn658);
V659:VNPU3_3 port map (start_vn,clk,rst,Lc659,C100V659,C479V659,C753V659,V659C100,V659C479,V659C753,SI659,end_vn659);
V660:VNPU3_3 port map (start_vn,clk,rst,Lc660,C101V660,C480V660,C754V660,V660C101,V660C480,V660C754,SI660,end_vn660);
V661:VNPU3_3 port map (start_vn,clk,rst,Lc661,C102V661,C385V661,C755V661,V661C102,V661C385,V661C755,SI661,end_vn661);
V662:VNPU3_3 port map (start_vn,clk,rst,Lc662,C103V662,C386V662,C756V662,V662C103,V662C386,V662C756,SI662,end_vn662);
V663:VNPU3_3 port map (start_vn,clk,rst,Lc663,C104V663,C387V663,C757V663,V663C104,V663C387,V663C757,SI663,end_vn663);
V664:VNPU3_3 port map (start_vn,clk,rst,Lc664,C105V664,C388V664,C758V664,V664C105,V664C388,V664C758,SI664,end_vn664);
V665:VNPU3_3 port map (start_vn,clk,rst,Lc665,C106V665,C389V665,C759V665,V665C106,V665C389,V665C759,SI665,end_vn665);
V666:VNPU3_3 port map (start_vn,clk,rst,Lc666,C107V666,C390V666,C760V666,V666C107,V666C390,V666C760,SI666,end_vn666);
V667:VNPU3_3 port map (start_vn,clk,rst,Lc667,C108V667,C391V667,C761V667,V667C108,V667C391,V667C761,SI667,end_vn667);
V668:VNPU3_3 port map (start_vn,clk,rst,Lc668,C109V668,C392V668,C762V668,V668C109,V668C392,V668C762,SI668,end_vn668);
V669:VNPU3_3 port map (start_vn,clk,rst,Lc669,C110V669,C393V669,C763V669,V669C110,V669C393,V669C763,SI669,end_vn669);
V670:VNPU3_3 port map (start_vn,clk,rst,Lc670,C111V670,C394V670,C764V670,V670C111,V670C394,V670C764,SI670,end_vn670);
V671:VNPU3_3 port map (start_vn,clk,rst,Lc671,C112V671,C395V671,C765V671,V671C112,V671C395,V671C765,SI671,end_vn671);
V672:VNPU3_3 port map (start_vn,clk,rst,Lc672,C113V672,C396V672,C766V672,V672C113,V672C396,V672C766,SI672,end_vn672);
V673:VNPU6_6 port map (start_vn,clk,rst,Lc673,C184V673,C256V673,C495V673,C822V673,C902V673,C1112V673,V673C184,V673C256,V673C495,V673C822,V673C902,V673C1112,SI673,end_vn673);
V674:VNPU6_6 port map (start_vn,clk,rst,Lc674,C185V674,C257V674,C496V674,C823V674,C903V674,C1113V674,V674C185,V674C257,V674C496,V674C823,V674C903,V674C1113,SI674,end_vn674);
V675:VNPU6_6 port map (start_vn,clk,rst,Lc675,C186V675,C258V675,C497V675,C824V675,C904V675,C1114V675,V675C186,V675C258,V675C497,V675C824,V675C904,V675C1114,SI675,end_vn675);
V676:VNPU6_6 port map (start_vn,clk,rst,Lc676,C187V676,C259V676,C498V676,C825V676,C905V676,C1115V676,V676C187,V676C259,V676C498,V676C825,V676C905,V676C1115,SI676,end_vn676);
V677:VNPU6_6 port map (start_vn,clk,rst,Lc677,C188V677,C260V677,C499V677,C826V677,C906V677,C1116V677,V677C188,V677C260,V677C499,V677C826,V677C906,V677C1116,SI677,end_vn677);
V678:VNPU6_6 port map (start_vn,clk,rst,Lc678,C189V678,C261V678,C500V678,C827V678,C907V678,C1117V678,V678C189,V678C261,V678C500,V678C827,V678C907,V678C1117,SI678,end_vn678);
V679:VNPU6_6 port map (start_vn,clk,rst,Lc679,C190V679,C262V679,C501V679,C828V679,C908V679,C1118V679,V679C190,V679C262,V679C501,V679C828,V679C908,V679C1118,SI679,end_vn679);
V680:VNPU6_6 port map (start_vn,clk,rst,Lc680,C191V680,C263V680,C502V680,C829V680,C909V680,C1119V680,V680C191,V680C263,V680C502,V680C829,V680C909,V680C1119,SI680,end_vn680);
V681:VNPU6_6 port map (start_vn,clk,rst,Lc681,C192V681,C264V681,C503V681,C830V681,C910V681,C1120V681,V681C192,V681C264,V681C503,V681C830,V681C910,V681C1120,SI681,end_vn681);
V682:VNPU6_6 port map (start_vn,clk,rst,Lc682,C97V682,C265V682,C504V682,C831V682,C911V682,C1121V682,V682C97,V682C265,V682C504,V682C831,V682C911,V682C1121,SI682,end_vn682);
V683:VNPU6_6 port map (start_vn,clk,rst,Lc683,C98V683,C266V683,C505V683,C832V683,C912V683,C1122V683,V683C98,V683C266,V683C505,V683C832,V683C912,V683C1122,SI683,end_vn683);
V684:VNPU6_6 port map (start_vn,clk,rst,Lc684,C99V684,C267V684,C506V684,C833V684,C913V684,C1123V684,V684C99,V684C267,V684C506,V684C833,V684C913,V684C1123,SI684,end_vn684);
V685:VNPU6_6 port map (start_vn,clk,rst,Lc685,C100V685,C268V685,C507V685,C834V685,C914V685,C1124V685,V685C100,V685C268,V685C507,V685C834,V685C914,V685C1124,SI685,end_vn685);
V686:VNPU6_6 port map (start_vn,clk,rst,Lc686,C101V686,C269V686,C508V686,C835V686,C915V686,C1125V686,V686C101,V686C269,V686C508,V686C835,V686C915,V686C1125,SI686,end_vn686);
V687:VNPU6_6 port map (start_vn,clk,rst,Lc687,C102V687,C270V687,C509V687,C836V687,C916V687,C1126V687,V687C102,V687C270,V687C509,V687C836,V687C916,V687C1126,SI687,end_vn687);
V688:VNPU6_6 port map (start_vn,clk,rst,Lc688,C103V688,C271V688,C510V688,C837V688,C917V688,C1127V688,V688C103,V688C271,V688C510,V688C837,V688C917,V688C1127,SI688,end_vn688);
V689:VNPU6_6 port map (start_vn,clk,rst,Lc689,C104V689,C272V689,C511V689,C838V689,C918V689,C1128V689,V689C104,V689C272,V689C511,V689C838,V689C918,V689C1128,SI689,end_vn689);
V690:VNPU6_6 port map (start_vn,clk,rst,Lc690,C105V690,C273V690,C512V690,C839V690,C919V690,C1129V690,V690C105,V690C273,V690C512,V690C839,V690C919,V690C1129,SI690,end_vn690);
V691:VNPU6_6 port map (start_vn,clk,rst,Lc691,C106V691,C274V691,C513V691,C840V691,C920V691,C1130V691,V691C106,V691C274,V691C513,V691C840,V691C920,V691C1130,SI691,end_vn691);
V692:VNPU6_6 port map (start_vn,clk,rst,Lc692,C107V692,C275V692,C514V692,C841V692,C921V692,C1131V692,V692C107,V692C275,V692C514,V692C841,V692C921,V692C1131,SI692,end_vn692);
V693:VNPU6_6 port map (start_vn,clk,rst,Lc693,C108V693,C276V693,C515V693,C842V693,C922V693,C1132V693,V693C108,V693C276,V693C515,V693C842,V693C922,V693C1132,SI693,end_vn693);
V694:VNPU6_6 port map (start_vn,clk,rst,Lc694,C109V694,C277V694,C516V694,C843V694,C923V694,C1133V694,V694C109,V694C277,V694C516,V694C843,V694C923,V694C1133,SI694,end_vn694);
V695:VNPU6_6 port map (start_vn,clk,rst,Lc695,C110V695,C278V695,C517V695,C844V695,C924V695,C1134V695,V695C110,V695C278,V695C517,V695C844,V695C924,V695C1134,SI695,end_vn695);
V696:VNPU6_6 port map (start_vn,clk,rst,Lc696,C111V696,C279V696,C518V696,C845V696,C925V696,C1135V696,V696C111,V696C279,V696C518,V696C845,V696C925,V696C1135,SI696,end_vn696);
V697:VNPU6_6 port map (start_vn,clk,rst,Lc697,C112V697,C280V697,C519V697,C846V697,C926V697,C1136V697,V697C112,V697C280,V697C519,V697C846,V697C926,V697C1136,SI697,end_vn697);
V698:VNPU6_6 port map (start_vn,clk,rst,Lc698,C113V698,C281V698,C520V698,C847V698,C927V698,C1137V698,V698C113,V698C281,V698C520,V698C847,V698C927,V698C1137,SI698,end_vn698);
V699:VNPU6_6 port map (start_vn,clk,rst,Lc699,C114V699,C282V699,C521V699,C848V699,C928V699,C1138V699,V699C114,V699C282,V699C521,V699C848,V699C928,V699C1138,SI699,end_vn699);
V700:VNPU6_6 port map (start_vn,clk,rst,Lc700,C115V700,C283V700,C522V700,C849V700,C929V700,C1139V700,V700C115,V700C283,V700C522,V700C849,V700C929,V700C1139,SI700,end_vn700);
V701:VNPU6_6 port map (start_vn,clk,rst,Lc701,C116V701,C284V701,C523V701,C850V701,C930V701,C1140V701,V701C116,V701C284,V701C523,V701C850,V701C930,V701C1140,SI701,end_vn701);
V702:VNPU6_6 port map (start_vn,clk,rst,Lc702,C117V702,C285V702,C524V702,C851V702,C931V702,C1141V702,V702C117,V702C285,V702C524,V702C851,V702C931,V702C1141,SI702,end_vn702);
V703:VNPU6_6 port map (start_vn,clk,rst,Lc703,C118V703,C286V703,C525V703,C852V703,C932V703,C1142V703,V703C118,V703C286,V703C525,V703C852,V703C932,V703C1142,SI703,end_vn703);
V704:VNPU6_6 port map (start_vn,clk,rst,Lc704,C119V704,C287V704,C526V704,C853V704,C933V704,C1143V704,V704C119,V704C287,V704C526,V704C853,V704C933,V704C1143,SI704,end_vn704);
V705:VNPU6_6 port map (start_vn,clk,rst,Lc705,C120V705,C288V705,C527V705,C854V705,C934V705,C1144V705,V705C120,V705C288,V705C527,V705C854,V705C934,V705C1144,SI705,end_vn705);
V706:VNPU6_6 port map (start_vn,clk,rst,Lc706,C121V706,C193V706,C528V706,C855V706,C935V706,C1145V706,V706C121,V706C193,V706C528,V706C855,V706C935,V706C1145,SI706,end_vn706);
V707:VNPU6_6 port map (start_vn,clk,rst,Lc707,C122V707,C194V707,C529V707,C856V707,C936V707,C1146V707,V707C122,V707C194,V707C529,V707C856,V707C936,V707C1146,SI707,end_vn707);
V708:VNPU6_6 port map (start_vn,clk,rst,Lc708,C123V708,C195V708,C530V708,C857V708,C937V708,C1147V708,V708C123,V708C195,V708C530,V708C857,V708C937,V708C1147,SI708,end_vn708);
V709:VNPU6_6 port map (start_vn,clk,rst,Lc709,C124V709,C196V709,C531V709,C858V709,C938V709,C1148V709,V709C124,V709C196,V709C531,V709C858,V709C938,V709C1148,SI709,end_vn709);
V710:VNPU6_6 port map (start_vn,clk,rst,Lc710,C125V710,C197V710,C532V710,C859V710,C939V710,C1149V710,V710C125,V710C197,V710C532,V710C859,V710C939,V710C1149,SI710,end_vn710);
V711:VNPU6_6 port map (start_vn,clk,rst,Lc711,C126V711,C198V711,C533V711,C860V711,C940V711,C1150V711,V711C126,V711C198,V711C533,V711C860,V711C940,V711C1150,SI711,end_vn711);
V712:VNPU6_6 port map (start_vn,clk,rst,Lc712,C127V712,C199V712,C534V712,C861V712,C941V712,C1151V712,V712C127,V712C199,V712C534,V712C861,V712C941,V712C1151,SI712,end_vn712);
V713:VNPU6_6 port map (start_vn,clk,rst,Lc713,C128V713,C200V713,C535V713,C862V713,C942V713,C1152V713,V713C128,V713C200,V713C535,V713C862,V713C942,V713C1152,SI713,end_vn713);
V714:VNPU6_6 port map (start_vn,clk,rst,Lc714,C129V714,C201V714,C536V714,C863V714,C943V714,C1057V714,V714C129,V714C201,V714C536,V714C863,V714C943,V714C1057,SI714,end_vn714);
V715:VNPU6_6 port map (start_vn,clk,rst,Lc715,C130V715,C202V715,C537V715,C864V715,C944V715,C1058V715,V715C130,V715C202,V715C537,V715C864,V715C944,V715C1058,SI715,end_vn715);
V716:VNPU6_6 port map (start_vn,clk,rst,Lc716,C131V716,C203V716,C538V716,C769V716,C945V716,C1059V716,V716C131,V716C203,V716C538,V716C769,V716C945,V716C1059,SI716,end_vn716);
V717:VNPU6_6 port map (start_vn,clk,rst,Lc717,C132V717,C204V717,C539V717,C770V717,C946V717,C1060V717,V717C132,V717C204,V717C539,V717C770,V717C946,V717C1060,SI717,end_vn717);
V718:VNPU6_6 port map (start_vn,clk,rst,Lc718,C133V718,C205V718,C540V718,C771V718,C947V718,C1061V718,V718C133,V718C205,V718C540,V718C771,V718C947,V718C1061,SI718,end_vn718);
V719:VNPU6_6 port map (start_vn,clk,rst,Lc719,C134V719,C206V719,C541V719,C772V719,C948V719,C1062V719,V719C134,V719C206,V719C541,V719C772,V719C948,V719C1062,SI719,end_vn719);
V720:VNPU6_6 port map (start_vn,clk,rst,Lc720,C135V720,C207V720,C542V720,C773V720,C949V720,C1063V720,V720C135,V720C207,V720C542,V720C773,V720C949,V720C1063,SI720,end_vn720);
V721:VNPU6_6 port map (start_vn,clk,rst,Lc721,C136V721,C208V721,C543V721,C774V721,C950V721,C1064V721,V721C136,V721C208,V721C543,V721C774,V721C950,V721C1064,SI721,end_vn721);
V722:VNPU6_6 port map (start_vn,clk,rst,Lc722,C137V722,C209V722,C544V722,C775V722,C951V722,C1065V722,V722C137,V722C209,V722C544,V722C775,V722C951,V722C1065,SI722,end_vn722);
V723:VNPU6_6 port map (start_vn,clk,rst,Lc723,C138V723,C210V723,C545V723,C776V723,C952V723,C1066V723,V723C138,V723C210,V723C545,V723C776,V723C952,V723C1066,SI723,end_vn723);
V724:VNPU6_6 port map (start_vn,clk,rst,Lc724,C139V724,C211V724,C546V724,C777V724,C953V724,C1067V724,V724C139,V724C211,V724C546,V724C777,V724C953,V724C1067,SI724,end_vn724);
V725:VNPU6_6 port map (start_vn,clk,rst,Lc725,C140V725,C212V725,C547V725,C778V725,C954V725,C1068V725,V725C140,V725C212,V725C547,V725C778,V725C954,V725C1068,SI725,end_vn725);
V726:VNPU6_6 port map (start_vn,clk,rst,Lc726,C141V726,C213V726,C548V726,C779V726,C955V726,C1069V726,V726C141,V726C213,V726C548,V726C779,V726C955,V726C1069,SI726,end_vn726);
V727:VNPU6_6 port map (start_vn,clk,rst,Lc727,C142V727,C214V727,C549V727,C780V727,C956V727,C1070V727,V727C142,V727C214,V727C549,V727C780,V727C956,V727C1070,SI727,end_vn727);
V728:VNPU6_6 port map (start_vn,clk,rst,Lc728,C143V728,C215V728,C550V728,C781V728,C957V728,C1071V728,V728C143,V728C215,V728C550,V728C781,V728C957,V728C1071,SI728,end_vn728);
V729:VNPU6_6 port map (start_vn,clk,rst,Lc729,C144V729,C216V729,C551V729,C782V729,C958V729,C1072V729,V729C144,V729C216,V729C551,V729C782,V729C958,V729C1072,SI729,end_vn729);
V730:VNPU6_6 port map (start_vn,clk,rst,Lc730,C145V730,C217V730,C552V730,C783V730,C959V730,C1073V730,V730C145,V730C217,V730C552,V730C783,V730C959,V730C1073,SI730,end_vn730);
V731:VNPU6_6 port map (start_vn,clk,rst,Lc731,C146V731,C218V731,C553V731,C784V731,C960V731,C1074V731,V731C146,V731C218,V731C553,V731C784,V731C960,V731C1074,SI731,end_vn731);
V732:VNPU6_6 port map (start_vn,clk,rst,Lc732,C147V732,C219V732,C554V732,C785V732,C865V732,C1075V732,V732C147,V732C219,V732C554,V732C785,V732C865,V732C1075,SI732,end_vn732);
V733:VNPU6_6 port map (start_vn,clk,rst,Lc733,C148V733,C220V733,C555V733,C786V733,C866V733,C1076V733,V733C148,V733C220,V733C555,V733C786,V733C866,V733C1076,SI733,end_vn733);
V734:VNPU6_6 port map (start_vn,clk,rst,Lc734,C149V734,C221V734,C556V734,C787V734,C867V734,C1077V734,V734C149,V734C221,V734C556,V734C787,V734C867,V734C1077,SI734,end_vn734);
V735:VNPU6_6 port map (start_vn,clk,rst,Lc735,C150V735,C222V735,C557V735,C788V735,C868V735,C1078V735,V735C150,V735C222,V735C557,V735C788,V735C868,V735C1078,SI735,end_vn735);
V736:VNPU6_6 port map (start_vn,clk,rst,Lc736,C151V736,C223V736,C558V736,C789V736,C869V736,C1079V736,V736C151,V736C223,V736C558,V736C789,V736C869,V736C1079,SI736,end_vn736);
V737:VNPU6_6 port map (start_vn,clk,rst,Lc737,C152V737,C224V737,C559V737,C790V737,C870V737,C1080V737,V737C152,V737C224,V737C559,V737C790,V737C870,V737C1080,SI737,end_vn737);
V738:VNPU6_6 port map (start_vn,clk,rst,Lc738,C153V738,C225V738,C560V738,C791V738,C871V738,C1081V738,V738C153,V738C225,V738C560,V738C791,V738C871,V738C1081,SI738,end_vn738);
V739:VNPU6_6 port map (start_vn,clk,rst,Lc739,C154V739,C226V739,C561V739,C792V739,C872V739,C1082V739,V739C154,V739C226,V739C561,V739C792,V739C872,V739C1082,SI739,end_vn739);
V740:VNPU6_6 port map (start_vn,clk,rst,Lc740,C155V740,C227V740,C562V740,C793V740,C873V740,C1083V740,V740C155,V740C227,V740C562,V740C793,V740C873,V740C1083,SI740,end_vn740);
V741:VNPU6_6 port map (start_vn,clk,rst,Lc741,C156V741,C228V741,C563V741,C794V741,C874V741,C1084V741,V741C156,V741C228,V741C563,V741C794,V741C874,V741C1084,SI741,end_vn741);
V742:VNPU6_6 port map (start_vn,clk,rst,Lc742,C157V742,C229V742,C564V742,C795V742,C875V742,C1085V742,V742C157,V742C229,V742C564,V742C795,V742C875,V742C1085,SI742,end_vn742);
V743:VNPU6_6 port map (start_vn,clk,rst,Lc743,C158V743,C230V743,C565V743,C796V743,C876V743,C1086V743,V743C158,V743C230,V743C565,V743C796,V743C876,V743C1086,SI743,end_vn743);
V744:VNPU6_6 port map (start_vn,clk,rst,Lc744,C159V744,C231V744,C566V744,C797V744,C877V744,C1087V744,V744C159,V744C231,V744C566,V744C797,V744C877,V744C1087,SI744,end_vn744);
V745:VNPU6_6 port map (start_vn,clk,rst,Lc745,C160V745,C232V745,C567V745,C798V745,C878V745,C1088V745,V745C160,V745C232,V745C567,V745C798,V745C878,V745C1088,SI745,end_vn745);
V746:VNPU6_6 port map (start_vn,clk,rst,Lc746,C161V746,C233V746,C568V746,C799V746,C879V746,C1089V746,V746C161,V746C233,V746C568,V746C799,V746C879,V746C1089,SI746,end_vn746);
V747:VNPU6_6 port map (start_vn,clk,rst,Lc747,C162V747,C234V747,C569V747,C800V747,C880V747,C1090V747,V747C162,V747C234,V747C569,V747C800,V747C880,V747C1090,SI747,end_vn747);
V748:VNPU6_6 port map (start_vn,clk,rst,Lc748,C163V748,C235V748,C570V748,C801V748,C881V748,C1091V748,V748C163,V748C235,V748C570,V748C801,V748C881,V748C1091,SI748,end_vn748);
V749:VNPU6_6 port map (start_vn,clk,rst,Lc749,C164V749,C236V749,C571V749,C802V749,C882V749,C1092V749,V749C164,V749C236,V749C571,V749C802,V749C882,V749C1092,SI749,end_vn749);
V750:VNPU6_6 port map (start_vn,clk,rst,Lc750,C165V750,C237V750,C572V750,C803V750,C883V750,C1093V750,V750C165,V750C237,V750C572,V750C803,V750C883,V750C1093,SI750,end_vn750);
V751:VNPU6_6 port map (start_vn,clk,rst,Lc751,C166V751,C238V751,C573V751,C804V751,C884V751,C1094V751,V751C166,V751C238,V751C573,V751C804,V751C884,V751C1094,SI751,end_vn751);
V752:VNPU6_6 port map (start_vn,clk,rst,Lc752,C167V752,C239V752,C574V752,C805V752,C885V752,C1095V752,V752C167,V752C239,V752C574,V752C805,V752C885,V752C1095,SI752,end_vn752);
V753:VNPU6_6 port map (start_vn,clk,rst,Lc753,C168V753,C240V753,C575V753,C806V753,C886V753,C1096V753,V753C168,V753C240,V753C575,V753C806,V753C886,V753C1096,SI753,end_vn753);
V754:VNPU6_6 port map (start_vn,clk,rst,Lc754,C169V754,C241V754,C576V754,C807V754,C887V754,C1097V754,V754C169,V754C241,V754C576,V754C807,V754C887,V754C1097,SI754,end_vn754);
V755:VNPU6_6 port map (start_vn,clk,rst,Lc755,C170V755,C242V755,C481V755,C808V755,C888V755,C1098V755,V755C170,V755C242,V755C481,V755C808,V755C888,V755C1098,SI755,end_vn755);
V756:VNPU6_6 port map (start_vn,clk,rst,Lc756,C171V756,C243V756,C482V756,C809V756,C889V756,C1099V756,V756C171,V756C243,V756C482,V756C809,V756C889,V756C1099,SI756,end_vn756);
V757:VNPU6_6 port map (start_vn,clk,rst,Lc757,C172V757,C244V757,C483V757,C810V757,C890V757,C1100V757,V757C172,V757C244,V757C483,V757C810,V757C890,V757C1100,SI757,end_vn757);
V758:VNPU6_6 port map (start_vn,clk,rst,Lc758,C173V758,C245V758,C484V758,C811V758,C891V758,C1101V758,V758C173,V758C245,V758C484,V758C811,V758C891,V758C1101,SI758,end_vn758);
V759:VNPU6_6 port map (start_vn,clk,rst,Lc759,C174V759,C246V759,C485V759,C812V759,C892V759,C1102V759,V759C174,V759C246,V759C485,V759C812,V759C892,V759C1102,SI759,end_vn759);
V760:VNPU6_6 port map (start_vn,clk,rst,Lc760,C175V760,C247V760,C486V760,C813V760,C893V760,C1103V760,V760C175,V760C247,V760C486,V760C813,V760C893,V760C1103,SI760,end_vn760);
V761:VNPU6_6 port map (start_vn,clk,rst,Lc761,C176V761,C248V761,C487V761,C814V761,C894V761,C1104V761,V761C176,V761C248,V761C487,V761C814,V761C894,V761C1104,SI761,end_vn761);
V762:VNPU6_6 port map (start_vn,clk,rst,Lc762,C177V762,C249V762,C488V762,C815V762,C895V762,C1105V762,V762C177,V762C249,V762C488,V762C815,V762C895,V762C1105,SI762,end_vn762);
V763:VNPU6_6 port map (start_vn,clk,rst,Lc763,C178V763,C250V763,C489V763,C816V763,C896V763,C1106V763,V763C178,V763C250,V763C489,V763C816,V763C896,V763C1106,SI763,end_vn763);
V764:VNPU6_6 port map (start_vn,clk,rst,Lc764,C179V764,C251V764,C490V764,C817V764,C897V764,C1107V764,V764C179,V764C251,V764C490,V764C817,V764C897,V764C1107,SI764,end_vn764);
V765:VNPU6_6 port map (start_vn,clk,rst,Lc765,C180V765,C252V765,C491V765,C818V765,C898V765,C1108V765,V765C180,V765C252,V765C491,V765C818,V765C898,V765C1108,SI765,end_vn765);
V766:VNPU6_6 port map (start_vn,clk,rst,Lc766,C181V766,C253V766,C492V766,C819V766,C899V766,C1109V766,V766C181,V766C253,V766C492,V766C819,V766C899,V766C1109,SI766,end_vn766);
V767:VNPU6_6 port map (start_vn,clk,rst,Lc767,C182V767,C254V767,C493V767,C820V767,C900V767,C1110V767,V767C182,V767C254,V767C493,V767C820,V767C900,V767C1110,SI767,end_vn767);
V768:VNPU6_6 port map (start_vn,clk,rst,Lc768,C183V768,C255V768,C494V768,C821V768,C901V768,C1111V768,V768C183,V768C255,V768C494,V768C821,V768C901,V768C1111,SI768,end_vn768);
V769:VNPU3_3 port map (start_vn,clk,rst,Lc769,C42V769,C320V769,C1018V769,V769C42,V769C320,V769C1018,SI769,end_vn769);
V770:VNPU3_3 port map (start_vn,clk,rst,Lc770,C43V770,C321V770,C1019V770,V770C43,V770C321,V770C1019,SI770,end_vn770);
V771:VNPU3_3 port map (start_vn,clk,rst,Lc771,C44V771,C322V771,C1020V771,V771C44,V771C322,V771C1020,SI771,end_vn771);
V772:VNPU3_3 port map (start_vn,clk,rst,Lc772,C45V772,C323V772,C1021V772,V772C45,V772C323,V772C1021,SI772,end_vn772);
V773:VNPU3_3 port map (start_vn,clk,rst,Lc773,C46V773,C324V773,C1022V773,V773C46,V773C324,V773C1022,SI773,end_vn773);
V774:VNPU3_3 port map (start_vn,clk,rst,Lc774,C47V774,C325V774,C1023V774,V774C47,V774C325,V774C1023,SI774,end_vn774);
V775:VNPU3_3 port map (start_vn,clk,rst,Lc775,C48V775,C326V775,C1024V775,V775C48,V775C326,V775C1024,SI775,end_vn775);
V776:VNPU3_3 port map (start_vn,clk,rst,Lc776,C49V776,C327V776,C1025V776,V776C49,V776C327,V776C1025,SI776,end_vn776);
V777:VNPU3_3 port map (start_vn,clk,rst,Lc777,C50V777,C328V777,C1026V777,V777C50,V777C328,V777C1026,SI777,end_vn777);
V778:VNPU3_3 port map (start_vn,clk,rst,Lc778,C51V778,C329V778,C1027V778,V778C51,V778C329,V778C1027,SI778,end_vn778);
V779:VNPU3_3 port map (start_vn,clk,rst,Lc779,C52V779,C330V779,C1028V779,V779C52,V779C330,V779C1028,SI779,end_vn779);
V780:VNPU3_3 port map (start_vn,clk,rst,Lc780,C53V780,C331V780,C1029V780,V780C53,V780C331,V780C1029,SI780,end_vn780);
V781:VNPU3_3 port map (start_vn,clk,rst,Lc781,C54V781,C332V781,C1030V781,V781C54,V781C332,V781C1030,SI781,end_vn781);
V782:VNPU3_3 port map (start_vn,clk,rst,Lc782,C55V782,C333V782,C1031V782,V782C55,V782C333,V782C1031,SI782,end_vn782);
V783:VNPU3_3 port map (start_vn,clk,rst,Lc783,C56V783,C334V783,C1032V783,V783C56,V783C334,V783C1032,SI783,end_vn783);
V784:VNPU3_3 port map (start_vn,clk,rst,Lc784,C57V784,C335V784,C1033V784,V784C57,V784C335,V784C1033,SI784,end_vn784);
V785:VNPU3_3 port map (start_vn,clk,rst,Lc785,C58V785,C336V785,C1034V785,V785C58,V785C336,V785C1034,SI785,end_vn785);
V786:VNPU3_3 port map (start_vn,clk,rst,Lc786,C59V786,C337V786,C1035V786,V786C59,V786C337,V786C1035,SI786,end_vn786);
V787:VNPU3_3 port map (start_vn,clk,rst,Lc787,C60V787,C338V787,C1036V787,V787C60,V787C338,V787C1036,SI787,end_vn787);
V788:VNPU3_3 port map (start_vn,clk,rst,Lc788,C61V788,C339V788,C1037V788,V788C61,V788C339,V788C1037,SI788,end_vn788);
V789:VNPU3_3 port map (start_vn,clk,rst,Lc789,C62V789,C340V789,C1038V789,V789C62,V789C340,V789C1038,SI789,end_vn789);
V790:VNPU3_3 port map (start_vn,clk,rst,Lc790,C63V790,C341V790,C1039V790,V790C63,V790C341,V790C1039,SI790,end_vn790);
V791:VNPU3_3 port map (start_vn,clk,rst,Lc791,C64V791,C342V791,C1040V791,V791C64,V791C342,V791C1040,SI791,end_vn791);
V792:VNPU3_3 port map (start_vn,clk,rst,Lc792,C65V792,C343V792,C1041V792,V792C65,V792C343,V792C1041,SI792,end_vn792);
V793:VNPU3_3 port map (start_vn,clk,rst,Lc793,C66V793,C344V793,C1042V793,V793C66,V793C344,V793C1042,SI793,end_vn793);
V794:VNPU3_3 port map (start_vn,clk,rst,Lc794,C67V794,C345V794,C1043V794,V794C67,V794C345,V794C1043,SI794,end_vn794);
V795:VNPU3_3 port map (start_vn,clk,rst,Lc795,C68V795,C346V795,C1044V795,V795C68,V795C346,V795C1044,SI795,end_vn795);
V796:VNPU3_3 port map (start_vn,clk,rst,Lc796,C69V796,C347V796,C1045V796,V796C69,V796C347,V796C1045,SI796,end_vn796);
V797:VNPU3_3 port map (start_vn,clk,rst,Lc797,C70V797,C348V797,C1046V797,V797C70,V797C348,V797C1046,SI797,end_vn797);
V798:VNPU3_3 port map (start_vn,clk,rst,Lc798,C71V798,C349V798,C1047V798,V798C71,V798C349,V798C1047,SI798,end_vn798);
V799:VNPU3_3 port map (start_vn,clk,rst,Lc799,C72V799,C350V799,C1048V799,V799C72,V799C350,V799C1048,SI799,end_vn799);
V800:VNPU3_3 port map (start_vn,clk,rst,Lc800,C73V800,C351V800,C1049V800,V800C73,V800C351,V800C1049,SI800,end_vn800);
V801:VNPU3_3 port map (start_vn,clk,rst,Lc801,C74V801,C352V801,C1050V801,V801C74,V801C352,V801C1050,SI801,end_vn801);
V802:VNPU3_3 port map (start_vn,clk,rst,Lc802,C75V802,C353V802,C1051V802,V802C75,V802C353,V802C1051,SI802,end_vn802);
V803:VNPU3_3 port map (start_vn,clk,rst,Lc803,C76V803,C354V803,C1052V803,V803C76,V803C354,V803C1052,SI803,end_vn803);
V804:VNPU3_3 port map (start_vn,clk,rst,Lc804,C77V804,C355V804,C1053V804,V804C77,V804C355,V804C1053,SI804,end_vn804);
V805:VNPU3_3 port map (start_vn,clk,rst,Lc805,C78V805,C356V805,C1054V805,V805C78,V805C356,V805C1054,SI805,end_vn805);
V806:VNPU3_3 port map (start_vn,clk,rst,Lc806,C79V806,C357V806,C1055V806,V806C79,V806C357,V806C1055,SI806,end_vn806);
V807:VNPU3_3 port map (start_vn,clk,rst,Lc807,C80V807,C358V807,C1056V807,V807C80,V807C358,V807C1056,SI807,end_vn807);
V808:VNPU3_3 port map (start_vn,clk,rst,Lc808,C81V808,C359V808,C961V808,V808C81,V808C359,V808C961,SI808,end_vn808);
V809:VNPU3_3 port map (start_vn,clk,rst,Lc809,C82V809,C360V809,C962V809,V809C82,V809C360,V809C962,SI809,end_vn809);
V810:VNPU3_3 port map (start_vn,clk,rst,Lc810,C83V810,C361V810,C963V810,V810C83,V810C361,V810C963,SI810,end_vn810);
V811:VNPU3_3 port map (start_vn,clk,rst,Lc811,C84V811,C362V811,C964V811,V811C84,V811C362,V811C964,SI811,end_vn811);
V812:VNPU3_3 port map (start_vn,clk,rst,Lc812,C85V812,C363V812,C965V812,V812C85,V812C363,V812C965,SI812,end_vn812);
V813:VNPU3_3 port map (start_vn,clk,rst,Lc813,C86V813,C364V813,C966V813,V813C86,V813C364,V813C966,SI813,end_vn813);
V814:VNPU3_3 port map (start_vn,clk,rst,Lc814,C87V814,C365V814,C967V814,V814C87,V814C365,V814C967,SI814,end_vn814);
V815:VNPU3_3 port map (start_vn,clk,rst,Lc815,C88V815,C366V815,C968V815,V815C88,V815C366,V815C968,SI815,end_vn815);
V816:VNPU3_3 port map (start_vn,clk,rst,Lc816,C89V816,C367V816,C969V816,V816C89,V816C367,V816C969,SI816,end_vn816);
V817:VNPU3_3 port map (start_vn,clk,rst,Lc817,C90V817,C368V817,C970V817,V817C90,V817C368,V817C970,SI817,end_vn817);
V818:VNPU3_3 port map (start_vn,clk,rst,Lc818,C91V818,C369V818,C971V818,V818C91,V818C369,V818C971,SI818,end_vn818);
V819:VNPU3_3 port map (start_vn,clk,rst,Lc819,C92V819,C370V819,C972V819,V819C92,V819C370,V819C972,SI819,end_vn819);
V820:VNPU3_3 port map (start_vn,clk,rst,Lc820,C93V820,C371V820,C973V820,V820C93,V820C371,V820C973,SI820,end_vn820);
V821:VNPU3_3 port map (start_vn,clk,rst,Lc821,C94V821,C372V821,C974V821,V821C94,V821C372,V821C974,SI821,end_vn821);
V822:VNPU3_3 port map (start_vn,clk,rst,Lc822,C95V822,C373V822,C975V822,V822C95,V822C373,V822C975,SI822,end_vn822);
V823:VNPU3_3 port map (start_vn,clk,rst,Lc823,C96V823,C374V823,C976V823,V823C96,V823C374,V823C976,SI823,end_vn823);
V824:VNPU3_3 port map (start_vn,clk,rst,Lc824,C1V824,C375V824,C977V824,V824C1,V824C375,V824C977,SI824,end_vn824);
V825:VNPU3_3 port map (start_vn,clk,rst,Lc825,C2V825,C376V825,C978V825,V825C2,V825C376,V825C978,SI825,end_vn825);
V826:VNPU3_3 port map (start_vn,clk,rst,Lc826,C3V826,C377V826,C979V826,V826C3,V826C377,V826C979,SI826,end_vn826);
V827:VNPU3_3 port map (start_vn,clk,rst,Lc827,C4V827,C378V827,C980V827,V827C4,V827C378,V827C980,SI827,end_vn827);
V828:VNPU3_3 port map (start_vn,clk,rst,Lc828,C5V828,C379V828,C981V828,V828C5,V828C379,V828C981,SI828,end_vn828);
V829:VNPU3_3 port map (start_vn,clk,rst,Lc829,C6V829,C380V829,C982V829,V829C6,V829C380,V829C982,SI829,end_vn829);
V830:VNPU3_3 port map (start_vn,clk,rst,Lc830,C7V830,C381V830,C983V830,V830C7,V830C381,V830C983,SI830,end_vn830);
V831:VNPU3_3 port map (start_vn,clk,rst,Lc831,C8V831,C382V831,C984V831,V831C8,V831C382,V831C984,SI831,end_vn831);
V832:VNPU3_3 port map (start_vn,clk,rst,Lc832,C9V832,C383V832,C985V832,V832C9,V832C383,V832C985,SI832,end_vn832);
V833:VNPU3_3 port map (start_vn,clk,rst,Lc833,C10V833,C384V833,C986V833,V833C10,V833C384,V833C986,SI833,end_vn833);
V834:VNPU3_3 port map (start_vn,clk,rst,Lc834,C11V834,C289V834,C987V834,V834C11,V834C289,V834C987,SI834,end_vn834);
V835:VNPU3_3 port map (start_vn,clk,rst,Lc835,C12V835,C290V835,C988V835,V835C12,V835C290,V835C988,SI835,end_vn835);
V836:VNPU3_3 port map (start_vn,clk,rst,Lc836,C13V836,C291V836,C989V836,V836C13,V836C291,V836C989,SI836,end_vn836);
V837:VNPU3_3 port map (start_vn,clk,rst,Lc837,C14V837,C292V837,C990V837,V837C14,V837C292,V837C990,SI837,end_vn837);
V838:VNPU3_3 port map (start_vn,clk,rst,Lc838,C15V838,C293V838,C991V838,V838C15,V838C293,V838C991,SI838,end_vn838);
V839:VNPU3_3 port map (start_vn,clk,rst,Lc839,C16V839,C294V839,C992V839,V839C16,V839C294,V839C992,SI839,end_vn839);
V840:VNPU3_3 port map (start_vn,clk,rst,Lc840,C17V840,C295V840,C993V840,V840C17,V840C295,V840C993,SI840,end_vn840);
V841:VNPU3_3 port map (start_vn,clk,rst,Lc841,C18V841,C296V841,C994V841,V841C18,V841C296,V841C994,SI841,end_vn841);
V842:VNPU3_3 port map (start_vn,clk,rst,Lc842,C19V842,C297V842,C995V842,V842C19,V842C297,V842C995,SI842,end_vn842);
V843:VNPU3_3 port map (start_vn,clk,rst,Lc843,C20V843,C298V843,C996V843,V843C20,V843C298,V843C996,SI843,end_vn843);
V844:VNPU3_3 port map (start_vn,clk,rst,Lc844,C21V844,C299V844,C997V844,V844C21,V844C299,V844C997,SI844,end_vn844);
V845:VNPU3_3 port map (start_vn,clk,rst,Lc845,C22V845,C300V845,C998V845,V845C22,V845C300,V845C998,SI845,end_vn845);
V846:VNPU3_3 port map (start_vn,clk,rst,Lc846,C23V846,C301V846,C999V846,V846C23,V846C301,V846C999,SI846,end_vn846);
V847:VNPU3_3 port map (start_vn,clk,rst,Lc847,C24V847,C302V847,C1000V847,V847C24,V847C302,V847C1000,SI847,end_vn847);
V848:VNPU3_3 port map (start_vn,clk,rst,Lc848,C25V848,C303V848,C1001V848,V848C25,V848C303,V848C1001,SI848,end_vn848);
V849:VNPU3_3 port map (start_vn,clk,rst,Lc849,C26V849,C304V849,C1002V849,V849C26,V849C304,V849C1002,SI849,end_vn849);
V850:VNPU3_3 port map (start_vn,clk,rst,Lc850,C27V850,C305V850,C1003V850,V850C27,V850C305,V850C1003,SI850,end_vn850);
V851:VNPU3_3 port map (start_vn,clk,rst,Lc851,C28V851,C306V851,C1004V851,V851C28,V851C306,V851C1004,SI851,end_vn851);
V852:VNPU3_3 port map (start_vn,clk,rst,Lc852,C29V852,C307V852,C1005V852,V852C29,V852C307,V852C1005,SI852,end_vn852);
V853:VNPU3_3 port map (start_vn,clk,rst,Lc853,C30V853,C308V853,C1006V853,V853C30,V853C308,V853C1006,SI853,end_vn853);
V854:VNPU3_3 port map (start_vn,clk,rst,Lc854,C31V854,C309V854,C1007V854,V854C31,V854C309,V854C1007,SI854,end_vn854);
V855:VNPU3_3 port map (start_vn,clk,rst,Lc855,C32V855,C310V855,C1008V855,V855C32,V855C310,V855C1008,SI855,end_vn855);
V856:VNPU3_3 port map (start_vn,clk,rst,Lc856,C33V856,C311V856,C1009V856,V856C33,V856C311,V856C1009,SI856,end_vn856);
V857:VNPU3_3 port map (start_vn,clk,rst,Lc857,C34V857,C312V857,C1010V857,V857C34,V857C312,V857C1010,SI857,end_vn857);
V858:VNPU3_3 port map (start_vn,clk,rst,Lc858,C35V858,C313V858,C1011V858,V858C35,V858C313,V858C1011,SI858,end_vn858);
V859:VNPU3_3 port map (start_vn,clk,rst,Lc859,C36V859,C314V859,C1012V859,V859C36,V859C314,V859C1012,SI859,end_vn859);
V860:VNPU3_3 port map (start_vn,clk,rst,Lc860,C37V860,C315V860,C1013V860,V860C37,V860C315,V860C1013,SI860,end_vn860);
V861:VNPU3_3 port map (start_vn,clk,rst,Lc861,C38V861,C316V861,C1014V861,V861C38,V861C316,V861C1014,SI861,end_vn861);
V862:VNPU3_3 port map (start_vn,clk,rst,Lc862,C39V862,C317V862,C1015V862,V862C39,V862C317,V862C1015,SI862,end_vn862);
V863:VNPU3_3 port map (start_vn,clk,rst,Lc863,C40V863,C318V863,C1016V863,V863C40,V863C318,V863C1016,SI863,end_vn863);
V864:VNPU3_3 port map (start_vn,clk,rst,Lc864,C41V864,C319V864,C1017V864,V864C41,V864C319,V864C1017,SI864,end_vn864);
V865:VNPU6_6 port map (start_vn,clk,rst,Lc865,C14V865,C360V865,C440V865,C659V865,C722V865,C1008V865,V865C14,V865C360,V865C440,V865C659,V865C722,V865C1008,SI865,end_vn865);
V866:VNPU6_6 port map (start_vn,clk,rst,Lc866,C15V866,C361V866,C441V866,C660V866,C723V866,C1009V866,V866C15,V866C361,V866C441,V866C660,V866C723,V866C1009,SI866,end_vn866);
V867:VNPU6_6 port map (start_vn,clk,rst,Lc867,C16V867,C362V867,C442V867,C661V867,C724V867,C1010V867,V867C16,V867C362,V867C442,V867C661,V867C724,V867C1010,SI867,end_vn867);
V868:VNPU6_6 port map (start_vn,clk,rst,Lc868,C17V868,C363V868,C443V868,C662V868,C725V868,C1011V868,V868C17,V868C363,V868C443,V868C662,V868C725,V868C1011,SI868,end_vn868);
V869:VNPU6_6 port map (start_vn,clk,rst,Lc869,C18V869,C364V869,C444V869,C663V869,C726V869,C1012V869,V869C18,V869C364,V869C444,V869C663,V869C726,V869C1012,SI869,end_vn869);
V870:VNPU6_6 port map (start_vn,clk,rst,Lc870,C19V870,C365V870,C445V870,C664V870,C727V870,C1013V870,V870C19,V870C365,V870C445,V870C664,V870C727,V870C1013,SI870,end_vn870);
V871:VNPU6_6 port map (start_vn,clk,rst,Lc871,C20V871,C366V871,C446V871,C665V871,C728V871,C1014V871,V871C20,V871C366,V871C446,V871C665,V871C728,V871C1014,SI871,end_vn871);
V872:VNPU6_6 port map (start_vn,clk,rst,Lc872,C21V872,C367V872,C447V872,C666V872,C729V872,C1015V872,V872C21,V872C367,V872C447,V872C666,V872C729,V872C1015,SI872,end_vn872);
V873:VNPU6_6 port map (start_vn,clk,rst,Lc873,C22V873,C368V873,C448V873,C667V873,C730V873,C1016V873,V873C22,V873C368,V873C448,V873C667,V873C730,V873C1016,SI873,end_vn873);
V874:VNPU6_6 port map (start_vn,clk,rst,Lc874,C23V874,C369V874,C449V874,C668V874,C731V874,C1017V874,V874C23,V874C369,V874C449,V874C668,V874C731,V874C1017,SI874,end_vn874);
V875:VNPU6_6 port map (start_vn,clk,rst,Lc875,C24V875,C370V875,C450V875,C669V875,C732V875,C1018V875,V875C24,V875C370,V875C450,V875C669,V875C732,V875C1018,SI875,end_vn875);
V876:VNPU6_6 port map (start_vn,clk,rst,Lc876,C25V876,C371V876,C451V876,C670V876,C733V876,C1019V876,V876C25,V876C371,V876C451,V876C670,V876C733,V876C1019,SI876,end_vn876);
V877:VNPU6_6 port map (start_vn,clk,rst,Lc877,C26V877,C372V877,C452V877,C671V877,C734V877,C1020V877,V877C26,V877C372,V877C452,V877C671,V877C734,V877C1020,SI877,end_vn877);
V878:VNPU6_6 port map (start_vn,clk,rst,Lc878,C27V878,C373V878,C453V878,C672V878,C735V878,C1021V878,V878C27,V878C373,V878C453,V878C672,V878C735,V878C1021,SI878,end_vn878);
V879:VNPU6_6 port map (start_vn,clk,rst,Lc879,C28V879,C374V879,C454V879,C577V879,C736V879,C1022V879,V879C28,V879C374,V879C454,V879C577,V879C736,V879C1022,SI879,end_vn879);
V880:VNPU6_6 port map (start_vn,clk,rst,Lc880,C29V880,C375V880,C455V880,C578V880,C737V880,C1023V880,V880C29,V880C375,V880C455,V880C578,V880C737,V880C1023,SI880,end_vn880);
V881:VNPU6_6 port map (start_vn,clk,rst,Lc881,C30V881,C376V881,C456V881,C579V881,C738V881,C1024V881,V881C30,V881C376,V881C456,V881C579,V881C738,V881C1024,SI881,end_vn881);
V882:VNPU6_6 port map (start_vn,clk,rst,Lc882,C31V882,C377V882,C457V882,C580V882,C739V882,C1025V882,V882C31,V882C377,V882C457,V882C580,V882C739,V882C1025,SI882,end_vn882);
V883:VNPU6_6 port map (start_vn,clk,rst,Lc883,C32V883,C378V883,C458V883,C581V883,C740V883,C1026V883,V883C32,V883C378,V883C458,V883C581,V883C740,V883C1026,SI883,end_vn883);
V884:VNPU6_6 port map (start_vn,clk,rst,Lc884,C33V884,C379V884,C459V884,C582V884,C741V884,C1027V884,V884C33,V884C379,V884C459,V884C582,V884C741,V884C1027,SI884,end_vn884);
V885:VNPU6_6 port map (start_vn,clk,rst,Lc885,C34V885,C380V885,C460V885,C583V885,C742V885,C1028V885,V885C34,V885C380,V885C460,V885C583,V885C742,V885C1028,SI885,end_vn885);
V886:VNPU6_6 port map (start_vn,clk,rst,Lc886,C35V886,C381V886,C461V886,C584V886,C743V886,C1029V886,V886C35,V886C381,V886C461,V886C584,V886C743,V886C1029,SI886,end_vn886);
V887:VNPU6_6 port map (start_vn,clk,rst,Lc887,C36V887,C382V887,C462V887,C585V887,C744V887,C1030V887,V887C36,V887C382,V887C462,V887C585,V887C744,V887C1030,SI887,end_vn887);
V888:VNPU6_6 port map (start_vn,clk,rst,Lc888,C37V888,C383V888,C463V888,C586V888,C745V888,C1031V888,V888C37,V888C383,V888C463,V888C586,V888C745,V888C1031,SI888,end_vn888);
V889:VNPU6_6 port map (start_vn,clk,rst,Lc889,C38V889,C384V889,C464V889,C587V889,C746V889,C1032V889,V889C38,V889C384,V889C464,V889C587,V889C746,V889C1032,SI889,end_vn889);
V890:VNPU6_6 port map (start_vn,clk,rst,Lc890,C39V890,C289V890,C465V890,C588V890,C747V890,C1033V890,V890C39,V890C289,V890C465,V890C588,V890C747,V890C1033,SI890,end_vn890);
V891:VNPU6_6 port map (start_vn,clk,rst,Lc891,C40V891,C290V891,C466V891,C589V891,C748V891,C1034V891,V891C40,V891C290,V891C466,V891C589,V891C748,V891C1034,SI891,end_vn891);
V892:VNPU6_6 port map (start_vn,clk,rst,Lc892,C41V892,C291V892,C467V892,C590V892,C749V892,C1035V892,V892C41,V892C291,V892C467,V892C590,V892C749,V892C1035,SI892,end_vn892);
V893:VNPU6_6 port map (start_vn,clk,rst,Lc893,C42V893,C292V893,C468V893,C591V893,C750V893,C1036V893,V893C42,V893C292,V893C468,V893C591,V893C750,V893C1036,SI893,end_vn893);
V894:VNPU6_6 port map (start_vn,clk,rst,Lc894,C43V894,C293V894,C469V894,C592V894,C751V894,C1037V894,V894C43,V894C293,V894C469,V894C592,V894C751,V894C1037,SI894,end_vn894);
V895:VNPU6_6 port map (start_vn,clk,rst,Lc895,C44V895,C294V895,C470V895,C593V895,C752V895,C1038V895,V895C44,V895C294,V895C470,V895C593,V895C752,V895C1038,SI895,end_vn895);
V896:VNPU6_6 port map (start_vn,clk,rst,Lc896,C45V896,C295V896,C471V896,C594V896,C753V896,C1039V896,V896C45,V896C295,V896C471,V896C594,V896C753,V896C1039,SI896,end_vn896);
V897:VNPU6_6 port map (start_vn,clk,rst,Lc897,C46V897,C296V897,C472V897,C595V897,C754V897,C1040V897,V897C46,V897C296,V897C472,V897C595,V897C754,V897C1040,SI897,end_vn897);
V898:VNPU6_6 port map (start_vn,clk,rst,Lc898,C47V898,C297V898,C473V898,C596V898,C755V898,C1041V898,V898C47,V898C297,V898C473,V898C596,V898C755,V898C1041,SI898,end_vn898);
V899:VNPU6_6 port map (start_vn,clk,rst,Lc899,C48V899,C298V899,C474V899,C597V899,C756V899,C1042V899,V899C48,V899C298,V899C474,V899C597,V899C756,V899C1042,SI899,end_vn899);
V900:VNPU6_6 port map (start_vn,clk,rst,Lc900,C49V900,C299V900,C475V900,C598V900,C757V900,C1043V900,V900C49,V900C299,V900C475,V900C598,V900C757,V900C1043,SI900,end_vn900);
V901:VNPU6_6 port map (start_vn,clk,rst,Lc901,C50V901,C300V901,C476V901,C599V901,C758V901,C1044V901,V901C50,V901C300,V901C476,V901C599,V901C758,V901C1044,SI901,end_vn901);
V902:VNPU6_6 port map (start_vn,clk,rst,Lc902,C51V902,C301V902,C477V902,C600V902,C759V902,C1045V902,V902C51,V902C301,V902C477,V902C600,V902C759,V902C1045,SI902,end_vn902);
V903:VNPU6_6 port map (start_vn,clk,rst,Lc903,C52V903,C302V903,C478V903,C601V903,C760V903,C1046V903,V903C52,V903C302,V903C478,V903C601,V903C760,V903C1046,SI903,end_vn903);
V904:VNPU6_6 port map (start_vn,clk,rst,Lc904,C53V904,C303V904,C479V904,C602V904,C761V904,C1047V904,V904C53,V904C303,V904C479,V904C602,V904C761,V904C1047,SI904,end_vn904);
V905:VNPU6_6 port map (start_vn,clk,rst,Lc905,C54V905,C304V905,C480V905,C603V905,C762V905,C1048V905,V905C54,V905C304,V905C480,V905C603,V905C762,V905C1048,SI905,end_vn905);
V906:VNPU6_6 port map (start_vn,clk,rst,Lc906,C55V906,C305V906,C385V906,C604V906,C763V906,C1049V906,V906C55,V906C305,V906C385,V906C604,V906C763,V906C1049,SI906,end_vn906);
V907:VNPU6_6 port map (start_vn,clk,rst,Lc907,C56V907,C306V907,C386V907,C605V907,C764V907,C1050V907,V907C56,V907C306,V907C386,V907C605,V907C764,V907C1050,SI907,end_vn907);
V908:VNPU6_6 port map (start_vn,clk,rst,Lc908,C57V908,C307V908,C387V908,C606V908,C765V908,C1051V908,V908C57,V908C307,V908C387,V908C606,V908C765,V908C1051,SI908,end_vn908);
V909:VNPU6_6 port map (start_vn,clk,rst,Lc909,C58V909,C308V909,C388V909,C607V909,C766V909,C1052V909,V909C58,V909C308,V909C388,V909C607,V909C766,V909C1052,SI909,end_vn909);
V910:VNPU6_6 port map (start_vn,clk,rst,Lc910,C59V910,C309V910,C389V910,C608V910,C767V910,C1053V910,V910C59,V910C309,V910C389,V910C608,V910C767,V910C1053,SI910,end_vn910);
V911:VNPU6_6 port map (start_vn,clk,rst,Lc911,C60V911,C310V911,C390V911,C609V911,C768V911,C1054V911,V911C60,V911C310,V911C390,V911C609,V911C768,V911C1054,SI911,end_vn911);
V912:VNPU6_6 port map (start_vn,clk,rst,Lc912,C61V912,C311V912,C391V912,C610V912,C673V912,C1055V912,V912C61,V912C311,V912C391,V912C610,V912C673,V912C1055,SI912,end_vn912);
V913:VNPU6_6 port map (start_vn,clk,rst,Lc913,C62V913,C312V913,C392V913,C611V913,C674V913,C1056V913,V913C62,V913C312,V913C392,V913C611,V913C674,V913C1056,SI913,end_vn913);
V914:VNPU6_6 port map (start_vn,clk,rst,Lc914,C63V914,C313V914,C393V914,C612V914,C675V914,C961V914,V914C63,V914C313,V914C393,V914C612,V914C675,V914C961,SI914,end_vn914);
V915:VNPU6_6 port map (start_vn,clk,rst,Lc915,C64V915,C314V915,C394V915,C613V915,C676V915,C962V915,V915C64,V915C314,V915C394,V915C613,V915C676,V915C962,SI915,end_vn915);
V916:VNPU6_6 port map (start_vn,clk,rst,Lc916,C65V916,C315V916,C395V916,C614V916,C677V916,C963V916,V916C65,V916C315,V916C395,V916C614,V916C677,V916C963,SI916,end_vn916);
V917:VNPU6_6 port map (start_vn,clk,rst,Lc917,C66V917,C316V917,C396V917,C615V917,C678V917,C964V917,V917C66,V917C316,V917C396,V917C615,V917C678,V917C964,SI917,end_vn917);
V918:VNPU6_6 port map (start_vn,clk,rst,Lc918,C67V918,C317V918,C397V918,C616V918,C679V918,C965V918,V918C67,V918C317,V918C397,V918C616,V918C679,V918C965,SI918,end_vn918);
V919:VNPU6_6 port map (start_vn,clk,rst,Lc919,C68V919,C318V919,C398V919,C617V919,C680V919,C966V919,V919C68,V919C318,V919C398,V919C617,V919C680,V919C966,SI919,end_vn919);
V920:VNPU6_6 port map (start_vn,clk,rst,Lc920,C69V920,C319V920,C399V920,C618V920,C681V920,C967V920,V920C69,V920C319,V920C399,V920C618,V920C681,V920C967,SI920,end_vn920);
V921:VNPU6_6 port map (start_vn,clk,rst,Lc921,C70V921,C320V921,C400V921,C619V921,C682V921,C968V921,V921C70,V921C320,V921C400,V921C619,V921C682,V921C968,SI921,end_vn921);
V922:VNPU6_6 port map (start_vn,clk,rst,Lc922,C71V922,C321V922,C401V922,C620V922,C683V922,C969V922,V922C71,V922C321,V922C401,V922C620,V922C683,V922C969,SI922,end_vn922);
V923:VNPU6_6 port map (start_vn,clk,rst,Lc923,C72V923,C322V923,C402V923,C621V923,C684V923,C970V923,V923C72,V923C322,V923C402,V923C621,V923C684,V923C970,SI923,end_vn923);
V924:VNPU6_6 port map (start_vn,clk,rst,Lc924,C73V924,C323V924,C403V924,C622V924,C685V924,C971V924,V924C73,V924C323,V924C403,V924C622,V924C685,V924C971,SI924,end_vn924);
V925:VNPU6_6 port map (start_vn,clk,rst,Lc925,C74V925,C324V925,C404V925,C623V925,C686V925,C972V925,V925C74,V925C324,V925C404,V925C623,V925C686,V925C972,SI925,end_vn925);
V926:VNPU6_6 port map (start_vn,clk,rst,Lc926,C75V926,C325V926,C405V926,C624V926,C687V926,C973V926,V926C75,V926C325,V926C405,V926C624,V926C687,V926C973,SI926,end_vn926);
V927:VNPU6_6 port map (start_vn,clk,rst,Lc927,C76V927,C326V927,C406V927,C625V927,C688V927,C974V927,V927C76,V927C326,V927C406,V927C625,V927C688,V927C974,SI927,end_vn927);
V928:VNPU6_6 port map (start_vn,clk,rst,Lc928,C77V928,C327V928,C407V928,C626V928,C689V928,C975V928,V928C77,V928C327,V928C407,V928C626,V928C689,V928C975,SI928,end_vn928);
V929:VNPU6_6 port map (start_vn,clk,rst,Lc929,C78V929,C328V929,C408V929,C627V929,C690V929,C976V929,V929C78,V929C328,V929C408,V929C627,V929C690,V929C976,SI929,end_vn929);
V930:VNPU6_6 port map (start_vn,clk,rst,Lc930,C79V930,C329V930,C409V930,C628V930,C691V930,C977V930,V930C79,V930C329,V930C409,V930C628,V930C691,V930C977,SI930,end_vn930);
V931:VNPU6_6 port map (start_vn,clk,rst,Lc931,C80V931,C330V931,C410V931,C629V931,C692V931,C978V931,V931C80,V931C330,V931C410,V931C629,V931C692,V931C978,SI931,end_vn931);
V932:VNPU6_6 port map (start_vn,clk,rst,Lc932,C81V932,C331V932,C411V932,C630V932,C693V932,C979V932,V932C81,V932C331,V932C411,V932C630,V932C693,V932C979,SI932,end_vn932);
V933:VNPU6_6 port map (start_vn,clk,rst,Lc933,C82V933,C332V933,C412V933,C631V933,C694V933,C980V933,V933C82,V933C332,V933C412,V933C631,V933C694,V933C980,SI933,end_vn933);
V934:VNPU6_6 port map (start_vn,clk,rst,Lc934,C83V934,C333V934,C413V934,C632V934,C695V934,C981V934,V934C83,V934C333,V934C413,V934C632,V934C695,V934C981,SI934,end_vn934);
V935:VNPU6_6 port map (start_vn,clk,rst,Lc935,C84V935,C334V935,C414V935,C633V935,C696V935,C982V935,V935C84,V935C334,V935C414,V935C633,V935C696,V935C982,SI935,end_vn935);
V936:VNPU6_6 port map (start_vn,clk,rst,Lc936,C85V936,C335V936,C415V936,C634V936,C697V936,C983V936,V936C85,V936C335,V936C415,V936C634,V936C697,V936C983,SI936,end_vn936);
V937:VNPU6_6 port map (start_vn,clk,rst,Lc937,C86V937,C336V937,C416V937,C635V937,C698V937,C984V937,V937C86,V937C336,V937C416,V937C635,V937C698,V937C984,SI937,end_vn937);
V938:VNPU6_6 port map (start_vn,clk,rst,Lc938,C87V938,C337V938,C417V938,C636V938,C699V938,C985V938,V938C87,V938C337,V938C417,V938C636,V938C699,V938C985,SI938,end_vn938);
V939:VNPU6_6 port map (start_vn,clk,rst,Lc939,C88V939,C338V939,C418V939,C637V939,C700V939,C986V939,V939C88,V939C338,V939C418,V939C637,V939C700,V939C986,SI939,end_vn939);
V940:VNPU6_6 port map (start_vn,clk,rst,Lc940,C89V940,C339V940,C419V940,C638V940,C701V940,C987V940,V940C89,V940C339,V940C419,V940C638,V940C701,V940C987,SI940,end_vn940);
V941:VNPU6_6 port map (start_vn,clk,rst,Lc941,C90V941,C340V941,C420V941,C639V941,C702V941,C988V941,V941C90,V941C340,V941C420,V941C639,V941C702,V941C988,SI941,end_vn941);
V942:VNPU6_6 port map (start_vn,clk,rst,Lc942,C91V942,C341V942,C421V942,C640V942,C703V942,C989V942,V942C91,V942C341,V942C421,V942C640,V942C703,V942C989,SI942,end_vn942);
V943:VNPU6_6 port map (start_vn,clk,rst,Lc943,C92V943,C342V943,C422V943,C641V943,C704V943,C990V943,V943C92,V943C342,V943C422,V943C641,V943C704,V943C990,SI943,end_vn943);
V944:VNPU6_6 port map (start_vn,clk,rst,Lc944,C93V944,C343V944,C423V944,C642V944,C705V944,C991V944,V944C93,V944C343,V944C423,V944C642,V944C705,V944C991,SI944,end_vn944);
V945:VNPU6_6 port map (start_vn,clk,rst,Lc945,C94V945,C344V945,C424V945,C643V945,C706V945,C992V945,V945C94,V945C344,V945C424,V945C643,V945C706,V945C992,SI945,end_vn945);
V946:VNPU6_6 port map (start_vn,clk,rst,Lc946,C95V946,C345V946,C425V946,C644V946,C707V946,C993V946,V946C95,V946C345,V946C425,V946C644,V946C707,V946C993,SI946,end_vn946);
V947:VNPU6_6 port map (start_vn,clk,rst,Lc947,C96V947,C346V947,C426V947,C645V947,C708V947,C994V947,V947C96,V947C346,V947C426,V947C645,V947C708,V947C994,SI947,end_vn947);
V948:VNPU6_6 port map (start_vn,clk,rst,Lc948,C1V948,C347V948,C427V948,C646V948,C709V948,C995V948,V948C1,V948C347,V948C427,V948C646,V948C709,V948C995,SI948,end_vn948);
V949:VNPU6_6 port map (start_vn,clk,rst,Lc949,C2V949,C348V949,C428V949,C647V949,C710V949,C996V949,V949C2,V949C348,V949C428,V949C647,V949C710,V949C996,SI949,end_vn949);
V950:VNPU6_6 port map (start_vn,clk,rst,Lc950,C3V950,C349V950,C429V950,C648V950,C711V950,C997V950,V950C3,V950C349,V950C429,V950C648,V950C711,V950C997,SI950,end_vn950);
V951:VNPU6_6 port map (start_vn,clk,rst,Lc951,C4V951,C350V951,C430V951,C649V951,C712V951,C998V951,V951C4,V951C350,V951C430,V951C649,V951C712,V951C998,SI951,end_vn951);
V952:VNPU6_6 port map (start_vn,clk,rst,Lc952,C5V952,C351V952,C431V952,C650V952,C713V952,C999V952,V952C5,V952C351,V952C431,V952C650,V952C713,V952C999,SI952,end_vn952);
V953:VNPU6_6 port map (start_vn,clk,rst,Lc953,C6V953,C352V953,C432V953,C651V953,C714V953,C1000V953,V953C6,V953C352,V953C432,V953C651,V953C714,V953C1000,SI953,end_vn953);
V954:VNPU6_6 port map (start_vn,clk,rst,Lc954,C7V954,C353V954,C433V954,C652V954,C715V954,C1001V954,V954C7,V954C353,V954C433,V954C652,V954C715,V954C1001,SI954,end_vn954);
V955:VNPU6_6 port map (start_vn,clk,rst,Lc955,C8V955,C354V955,C434V955,C653V955,C716V955,C1002V955,V955C8,V955C354,V955C434,V955C653,V955C716,V955C1002,SI955,end_vn955);
V956:VNPU6_6 port map (start_vn,clk,rst,Lc956,C9V956,C355V956,C435V956,C654V956,C717V956,C1003V956,V956C9,V956C355,V956C435,V956C654,V956C717,V956C1003,SI956,end_vn956);
V957:VNPU6_6 port map (start_vn,clk,rst,Lc957,C10V957,C356V957,C436V957,C655V957,C718V957,C1004V957,V957C10,V957C356,V957C436,V957C655,V957C718,V957C1004,SI957,end_vn957);
V958:VNPU6_6 port map (start_vn,clk,rst,Lc958,C11V958,C357V958,C437V958,C656V958,C719V958,C1005V958,V958C11,V958C357,V958C437,V958C656,V958C719,V958C1005,SI958,end_vn958);
V959:VNPU6_6 port map (start_vn,clk,rst,Lc959,C12V959,C358V959,C438V959,C657V959,C720V959,C1006V959,V959C12,V959C358,V959C438,V959C657,V959C720,V959C1006,SI959,end_vn959);
V960:VNPU6_6 port map (start_vn,clk,rst,Lc960,C13V960,C359V960,C439V960,C658V960,C721V960,C1007V960,V960C13,V960C359,V960C439,V960C658,V960C721,V960C1007,SI960,end_vn960);
V961:VNPU3_3 port map (start_vn,clk,rst,Lc961,C409V961,C655V961,C891V961,V961C409,V961C655,V961C891,SI961,end_vn961);
V962:VNPU3_3 port map (start_vn,clk,rst,Lc962,C410V962,C656V962,C892V962,V962C410,V962C656,V962C892,SI962,end_vn962);
V963:VNPU3_3 port map (start_vn,clk,rst,Lc963,C411V963,C657V963,C893V963,V963C411,V963C657,V963C893,SI963,end_vn963);
V964:VNPU3_3 port map (start_vn,clk,rst,Lc964,C412V964,C658V964,C894V964,V964C412,V964C658,V964C894,SI964,end_vn964);
V965:VNPU3_3 port map (start_vn,clk,rst,Lc965,C413V965,C659V965,C895V965,V965C413,V965C659,V965C895,SI965,end_vn965);
V966:VNPU3_3 port map (start_vn,clk,rst,Lc966,C414V966,C660V966,C896V966,V966C414,V966C660,V966C896,SI966,end_vn966);
V967:VNPU3_3 port map (start_vn,clk,rst,Lc967,C415V967,C661V967,C897V967,V967C415,V967C661,V967C897,SI967,end_vn967);
V968:VNPU3_3 port map (start_vn,clk,rst,Lc968,C416V968,C662V968,C898V968,V968C416,V968C662,V968C898,SI968,end_vn968);
V969:VNPU3_3 port map (start_vn,clk,rst,Lc969,C417V969,C663V969,C899V969,V969C417,V969C663,V969C899,SI969,end_vn969);
V970:VNPU3_3 port map (start_vn,clk,rst,Lc970,C418V970,C664V970,C900V970,V970C418,V970C664,V970C900,SI970,end_vn970);
V971:VNPU3_3 port map (start_vn,clk,rst,Lc971,C419V971,C665V971,C901V971,V971C419,V971C665,V971C901,SI971,end_vn971);
V972:VNPU3_3 port map (start_vn,clk,rst,Lc972,C420V972,C666V972,C902V972,V972C420,V972C666,V972C902,SI972,end_vn972);
V973:VNPU3_3 port map (start_vn,clk,rst,Lc973,C421V973,C667V973,C903V973,V973C421,V973C667,V973C903,SI973,end_vn973);
V974:VNPU3_3 port map (start_vn,clk,rst,Lc974,C422V974,C668V974,C904V974,V974C422,V974C668,V974C904,SI974,end_vn974);
V975:VNPU3_3 port map (start_vn,clk,rst,Lc975,C423V975,C669V975,C905V975,V975C423,V975C669,V975C905,SI975,end_vn975);
V976:VNPU3_3 port map (start_vn,clk,rst,Lc976,C424V976,C670V976,C906V976,V976C424,V976C670,V976C906,SI976,end_vn976);
V977:VNPU3_3 port map (start_vn,clk,rst,Lc977,C425V977,C671V977,C907V977,V977C425,V977C671,V977C907,SI977,end_vn977);
V978:VNPU3_3 port map (start_vn,clk,rst,Lc978,C426V978,C672V978,C908V978,V978C426,V978C672,V978C908,SI978,end_vn978);
V979:VNPU3_3 port map (start_vn,clk,rst,Lc979,C427V979,C577V979,C909V979,V979C427,V979C577,V979C909,SI979,end_vn979);
V980:VNPU3_3 port map (start_vn,clk,rst,Lc980,C428V980,C578V980,C910V980,V980C428,V980C578,V980C910,SI980,end_vn980);
V981:VNPU3_3 port map (start_vn,clk,rst,Lc981,C429V981,C579V981,C911V981,V981C429,V981C579,V981C911,SI981,end_vn981);
V982:VNPU3_3 port map (start_vn,clk,rst,Lc982,C430V982,C580V982,C912V982,V982C430,V982C580,V982C912,SI982,end_vn982);
V983:VNPU3_3 port map (start_vn,clk,rst,Lc983,C431V983,C581V983,C913V983,V983C431,V983C581,V983C913,SI983,end_vn983);
V984:VNPU3_3 port map (start_vn,clk,rst,Lc984,C432V984,C582V984,C914V984,V984C432,V984C582,V984C914,SI984,end_vn984);
V985:VNPU3_3 port map (start_vn,clk,rst,Lc985,C433V985,C583V985,C915V985,V985C433,V985C583,V985C915,SI985,end_vn985);
V986:VNPU3_3 port map (start_vn,clk,rst,Lc986,C434V986,C584V986,C916V986,V986C434,V986C584,V986C916,SI986,end_vn986);
V987:VNPU3_3 port map (start_vn,clk,rst,Lc987,C435V987,C585V987,C917V987,V987C435,V987C585,V987C917,SI987,end_vn987);
V988:VNPU3_3 port map (start_vn,clk,rst,Lc988,C436V988,C586V988,C918V988,V988C436,V988C586,V988C918,SI988,end_vn988);
V989:VNPU3_3 port map (start_vn,clk,rst,Lc989,C437V989,C587V989,C919V989,V989C437,V989C587,V989C919,SI989,end_vn989);
V990:VNPU3_3 port map (start_vn,clk,rst,Lc990,C438V990,C588V990,C920V990,V990C438,V990C588,V990C920,SI990,end_vn990);
V991:VNPU3_3 port map (start_vn,clk,rst,Lc991,C439V991,C589V991,C921V991,V991C439,V991C589,V991C921,SI991,end_vn991);
V992:VNPU3_3 port map (start_vn,clk,rst,Lc992,C440V992,C590V992,C922V992,V992C440,V992C590,V992C922,SI992,end_vn992);
V993:VNPU3_3 port map (start_vn,clk,rst,Lc993,C441V993,C591V993,C923V993,V993C441,V993C591,V993C923,SI993,end_vn993);
V994:VNPU3_3 port map (start_vn,clk,rst,Lc994,C442V994,C592V994,C924V994,V994C442,V994C592,V994C924,SI994,end_vn994);
V995:VNPU3_3 port map (start_vn,clk,rst,Lc995,C443V995,C593V995,C925V995,V995C443,V995C593,V995C925,SI995,end_vn995);
V996:VNPU3_3 port map (start_vn,clk,rst,Lc996,C444V996,C594V996,C926V996,V996C444,V996C594,V996C926,SI996,end_vn996);
V997:VNPU3_3 port map (start_vn,clk,rst,Lc997,C445V997,C595V997,C927V997,V997C445,V997C595,V997C927,SI997,end_vn997);
V998:VNPU3_3 port map (start_vn,clk,rst,Lc998,C446V998,C596V998,C928V998,V998C446,V998C596,V998C928,SI998,end_vn998);
V999:VNPU3_3 port map (start_vn,clk,rst,Lc999,C447V999,C597V999,C929V999,V999C447,V999C597,V999C929,SI999,end_vn999);
V1000:VNPU3_3 port map (start_vn,clk,rst,Lc1000,C448V1000,C598V1000,C930V1000,V1000C448,V1000C598,V1000C930,SI1000,end_vn1000);
V1001:VNPU3_3 port map (start_vn,clk,rst,Lc1001,C449V1001,C599V1001,C931V1001,V1001C449,V1001C599,V1001C931,SI1001,end_vn1001);
V1002:VNPU3_3 port map (start_vn,clk,rst,Lc1002,C450V1002,C600V1002,C932V1002,V1002C450,V1002C600,V1002C932,SI1002,end_vn1002);
V1003:VNPU3_3 port map (start_vn,clk,rst,Lc1003,C451V1003,C601V1003,C933V1003,V1003C451,V1003C601,V1003C933,SI1003,end_vn1003);
V1004:VNPU3_3 port map (start_vn,clk,rst,Lc1004,C452V1004,C602V1004,C934V1004,V1004C452,V1004C602,V1004C934,SI1004,end_vn1004);
V1005:VNPU3_3 port map (start_vn,clk,rst,Lc1005,C453V1005,C603V1005,C935V1005,V1005C453,V1005C603,V1005C935,SI1005,end_vn1005);
V1006:VNPU3_3 port map (start_vn,clk,rst,Lc1006,C454V1006,C604V1006,C936V1006,V1006C454,V1006C604,V1006C936,SI1006,end_vn1006);
V1007:VNPU3_3 port map (start_vn,clk,rst,Lc1007,C455V1007,C605V1007,C937V1007,V1007C455,V1007C605,V1007C937,SI1007,end_vn1007);
V1008:VNPU3_3 port map (start_vn,clk,rst,Lc1008,C456V1008,C606V1008,C938V1008,V1008C456,V1008C606,V1008C938,SI1008,end_vn1008);
V1009:VNPU3_3 port map (start_vn,clk,rst,Lc1009,C457V1009,C607V1009,C939V1009,V1009C457,V1009C607,V1009C939,SI1009,end_vn1009);
V1010:VNPU3_3 port map (start_vn,clk,rst,Lc1010,C458V1010,C608V1010,C940V1010,V1010C458,V1010C608,V1010C940,SI1010,end_vn1010);
V1011:VNPU3_3 port map (start_vn,clk,rst,Lc1011,C459V1011,C609V1011,C941V1011,V1011C459,V1011C609,V1011C941,SI1011,end_vn1011);
V1012:VNPU3_3 port map (start_vn,clk,rst,Lc1012,C460V1012,C610V1012,C942V1012,V1012C460,V1012C610,V1012C942,SI1012,end_vn1012);
V1013:VNPU3_3 port map (start_vn,clk,rst,Lc1013,C461V1013,C611V1013,C943V1013,V1013C461,V1013C611,V1013C943,SI1013,end_vn1013);
V1014:VNPU3_3 port map (start_vn,clk,rst,Lc1014,C462V1014,C612V1014,C944V1014,V1014C462,V1014C612,V1014C944,SI1014,end_vn1014);
V1015:VNPU3_3 port map (start_vn,clk,rst,Lc1015,C463V1015,C613V1015,C945V1015,V1015C463,V1015C613,V1015C945,SI1015,end_vn1015);
V1016:VNPU3_3 port map (start_vn,clk,rst,Lc1016,C464V1016,C614V1016,C946V1016,V1016C464,V1016C614,V1016C946,SI1016,end_vn1016);
V1017:VNPU3_3 port map (start_vn,clk,rst,Lc1017,C465V1017,C615V1017,C947V1017,V1017C465,V1017C615,V1017C947,SI1017,end_vn1017);
V1018:VNPU3_3 port map (start_vn,clk,rst,Lc1018,C466V1018,C616V1018,C948V1018,V1018C466,V1018C616,V1018C948,SI1018,end_vn1018);
V1019:VNPU3_3 port map (start_vn,clk,rst,Lc1019,C467V1019,C617V1019,C949V1019,V1019C467,V1019C617,V1019C949,SI1019,end_vn1019);
V1020:VNPU3_3 port map (start_vn,clk,rst,Lc1020,C468V1020,C618V1020,C950V1020,V1020C468,V1020C618,V1020C950,SI1020,end_vn1020);
V1021:VNPU3_3 port map (start_vn,clk,rst,Lc1021,C469V1021,C619V1021,C951V1021,V1021C469,V1021C619,V1021C951,SI1021,end_vn1021);
V1022:VNPU3_3 port map (start_vn,clk,rst,Lc1022,C470V1022,C620V1022,C952V1022,V1022C470,V1022C620,V1022C952,SI1022,end_vn1022);
V1023:VNPU3_3 port map (start_vn,clk,rst,Lc1023,C471V1023,C621V1023,C953V1023,V1023C471,V1023C621,V1023C953,SI1023,end_vn1023);
V1024:VNPU3_3 port map (start_vn,clk,rst,Lc1024,C472V1024,C622V1024,C954V1024,V1024C472,V1024C622,V1024C954,SI1024,end_vn1024);
V1025:VNPU3_3 port map (start_vn,clk,rst,Lc1025,C473V1025,C623V1025,C955V1025,V1025C473,V1025C623,V1025C955,SI1025,end_vn1025);
V1026:VNPU3_3 port map (start_vn,clk,rst,Lc1026,C474V1026,C624V1026,C956V1026,V1026C474,V1026C624,V1026C956,SI1026,end_vn1026);
V1027:VNPU3_3 port map (start_vn,clk,rst,Lc1027,C475V1027,C625V1027,C957V1027,V1027C475,V1027C625,V1027C957,SI1027,end_vn1027);
V1028:VNPU3_3 port map (start_vn,clk,rst,Lc1028,C476V1028,C626V1028,C958V1028,V1028C476,V1028C626,V1028C958,SI1028,end_vn1028);
V1029:VNPU3_3 port map (start_vn,clk,rst,Lc1029,C477V1029,C627V1029,C959V1029,V1029C477,V1029C627,V1029C959,SI1029,end_vn1029);
V1030:VNPU3_3 port map (start_vn,clk,rst,Lc1030,C478V1030,C628V1030,C960V1030,V1030C478,V1030C628,V1030C960,SI1030,end_vn1030);
V1031:VNPU3_3 port map (start_vn,clk,rst,Lc1031,C479V1031,C629V1031,C865V1031,V1031C479,V1031C629,V1031C865,SI1031,end_vn1031);
V1032:VNPU3_3 port map (start_vn,clk,rst,Lc1032,C480V1032,C630V1032,C866V1032,V1032C480,V1032C630,V1032C866,SI1032,end_vn1032);
V1033:VNPU3_3 port map (start_vn,clk,rst,Lc1033,C385V1033,C631V1033,C867V1033,V1033C385,V1033C631,V1033C867,SI1033,end_vn1033);
V1034:VNPU3_3 port map (start_vn,clk,rst,Lc1034,C386V1034,C632V1034,C868V1034,V1034C386,V1034C632,V1034C868,SI1034,end_vn1034);
V1035:VNPU3_3 port map (start_vn,clk,rst,Lc1035,C387V1035,C633V1035,C869V1035,V1035C387,V1035C633,V1035C869,SI1035,end_vn1035);
V1036:VNPU3_3 port map (start_vn,clk,rst,Lc1036,C388V1036,C634V1036,C870V1036,V1036C388,V1036C634,V1036C870,SI1036,end_vn1036);
V1037:VNPU3_3 port map (start_vn,clk,rst,Lc1037,C389V1037,C635V1037,C871V1037,V1037C389,V1037C635,V1037C871,SI1037,end_vn1037);
V1038:VNPU3_3 port map (start_vn,clk,rst,Lc1038,C390V1038,C636V1038,C872V1038,V1038C390,V1038C636,V1038C872,SI1038,end_vn1038);
V1039:VNPU3_3 port map (start_vn,clk,rst,Lc1039,C391V1039,C637V1039,C873V1039,V1039C391,V1039C637,V1039C873,SI1039,end_vn1039);
V1040:VNPU3_3 port map (start_vn,clk,rst,Lc1040,C392V1040,C638V1040,C874V1040,V1040C392,V1040C638,V1040C874,SI1040,end_vn1040);
V1041:VNPU3_3 port map (start_vn,clk,rst,Lc1041,C393V1041,C639V1041,C875V1041,V1041C393,V1041C639,V1041C875,SI1041,end_vn1041);
V1042:VNPU3_3 port map (start_vn,clk,rst,Lc1042,C394V1042,C640V1042,C876V1042,V1042C394,V1042C640,V1042C876,SI1042,end_vn1042);
V1043:VNPU3_3 port map (start_vn,clk,rst,Lc1043,C395V1043,C641V1043,C877V1043,V1043C395,V1043C641,V1043C877,SI1043,end_vn1043);
V1044:VNPU3_3 port map (start_vn,clk,rst,Lc1044,C396V1044,C642V1044,C878V1044,V1044C396,V1044C642,V1044C878,SI1044,end_vn1044);
V1045:VNPU3_3 port map (start_vn,clk,rst,Lc1045,C397V1045,C643V1045,C879V1045,V1045C397,V1045C643,V1045C879,SI1045,end_vn1045);
V1046:VNPU3_3 port map (start_vn,clk,rst,Lc1046,C398V1046,C644V1046,C880V1046,V1046C398,V1046C644,V1046C880,SI1046,end_vn1046);
V1047:VNPU3_3 port map (start_vn,clk,rst,Lc1047,C399V1047,C645V1047,C881V1047,V1047C399,V1047C645,V1047C881,SI1047,end_vn1047);
V1048:VNPU3_3 port map (start_vn,clk,rst,Lc1048,C400V1048,C646V1048,C882V1048,V1048C400,V1048C646,V1048C882,SI1048,end_vn1048);
V1049:VNPU3_3 port map (start_vn,clk,rst,Lc1049,C401V1049,C647V1049,C883V1049,V1049C401,V1049C647,V1049C883,SI1049,end_vn1049);
V1050:VNPU3_3 port map (start_vn,clk,rst,Lc1050,C402V1050,C648V1050,C884V1050,V1050C402,V1050C648,V1050C884,SI1050,end_vn1050);
V1051:VNPU3_3 port map (start_vn,clk,rst,Lc1051,C403V1051,C649V1051,C885V1051,V1051C403,V1051C649,V1051C885,SI1051,end_vn1051);
V1052:VNPU3_3 port map (start_vn,clk,rst,Lc1052,C404V1052,C650V1052,C886V1052,V1052C404,V1052C650,V1052C886,SI1052,end_vn1052);
V1053:VNPU3_3 port map (start_vn,clk,rst,Lc1053,C405V1053,C651V1053,C887V1053,V1053C405,V1053C651,V1053C887,SI1053,end_vn1053);
V1054:VNPU3_3 port map (start_vn,clk,rst,Lc1054,C406V1054,C652V1054,C888V1054,V1054C406,V1054C652,V1054C888,SI1054,end_vn1054);
V1055:VNPU3_3 port map (start_vn,clk,rst,Lc1055,C407V1055,C653V1055,C889V1055,V1055C407,V1055C653,V1055C889,SI1055,end_vn1055);
V1056:VNPU3_3 port map (start_vn,clk,rst,Lc1056,C408V1056,C654V1056,C890V1056,V1056C408,V1056C654,V1056C890,SI1056,end_vn1056);
V1057:VNPU6_6 port map (start_vn,clk,rst,Lc1057,C181V1057,C193V1057,C498V1057,C814V1057,C889V1057,C1127V1057,V1057C181,V1057C193,V1057C498,V1057C814,V1057C889,V1057C1127,SI1057,end_vn1057);
V1058:VNPU6_6 port map (start_vn,clk,rst,Lc1058,C182V1058,C194V1058,C499V1058,C815V1058,C890V1058,C1128V1058,V1058C182,V1058C194,V1058C499,V1058C815,V1058C890,V1058C1128,SI1058,end_vn1058);
V1059:VNPU6_6 port map (start_vn,clk,rst,Lc1059,C183V1059,C195V1059,C500V1059,C816V1059,C891V1059,C1129V1059,V1059C183,V1059C195,V1059C500,V1059C816,V1059C891,V1059C1129,SI1059,end_vn1059);
V1060:VNPU6_6 port map (start_vn,clk,rst,Lc1060,C184V1060,C196V1060,C501V1060,C817V1060,C892V1060,C1130V1060,V1060C184,V1060C196,V1060C501,V1060C817,V1060C892,V1060C1130,SI1060,end_vn1060);
V1061:VNPU6_6 port map (start_vn,clk,rst,Lc1061,C185V1061,C197V1061,C502V1061,C818V1061,C893V1061,C1131V1061,V1061C185,V1061C197,V1061C502,V1061C818,V1061C893,V1061C1131,SI1061,end_vn1061);
V1062:VNPU6_6 port map (start_vn,clk,rst,Lc1062,C186V1062,C198V1062,C503V1062,C819V1062,C894V1062,C1132V1062,V1062C186,V1062C198,V1062C503,V1062C819,V1062C894,V1062C1132,SI1062,end_vn1062);
V1063:VNPU6_6 port map (start_vn,clk,rst,Lc1063,C187V1063,C199V1063,C504V1063,C820V1063,C895V1063,C1133V1063,V1063C187,V1063C199,V1063C504,V1063C820,V1063C895,V1063C1133,SI1063,end_vn1063);
V1064:VNPU6_6 port map (start_vn,clk,rst,Lc1064,C188V1064,C200V1064,C505V1064,C821V1064,C896V1064,C1134V1064,V1064C188,V1064C200,V1064C505,V1064C821,V1064C896,V1064C1134,SI1064,end_vn1064);
V1065:VNPU6_6 port map (start_vn,clk,rst,Lc1065,C189V1065,C201V1065,C506V1065,C822V1065,C897V1065,C1135V1065,V1065C189,V1065C201,V1065C506,V1065C822,V1065C897,V1065C1135,SI1065,end_vn1065);
V1066:VNPU6_6 port map (start_vn,clk,rst,Lc1066,C190V1066,C202V1066,C507V1066,C823V1066,C898V1066,C1136V1066,V1066C190,V1066C202,V1066C507,V1066C823,V1066C898,V1066C1136,SI1066,end_vn1066);
V1067:VNPU6_6 port map (start_vn,clk,rst,Lc1067,C191V1067,C203V1067,C508V1067,C824V1067,C899V1067,C1137V1067,V1067C191,V1067C203,V1067C508,V1067C824,V1067C899,V1067C1137,SI1067,end_vn1067);
V1068:VNPU6_6 port map (start_vn,clk,rst,Lc1068,C192V1068,C204V1068,C509V1068,C825V1068,C900V1068,C1138V1068,V1068C192,V1068C204,V1068C509,V1068C825,V1068C900,V1068C1138,SI1068,end_vn1068);
V1069:VNPU6_6 port map (start_vn,clk,rst,Lc1069,C97V1069,C205V1069,C510V1069,C826V1069,C901V1069,C1139V1069,V1069C97,V1069C205,V1069C510,V1069C826,V1069C901,V1069C1139,SI1069,end_vn1069);
V1070:VNPU6_6 port map (start_vn,clk,rst,Lc1070,C98V1070,C206V1070,C511V1070,C827V1070,C902V1070,C1140V1070,V1070C98,V1070C206,V1070C511,V1070C827,V1070C902,V1070C1140,SI1070,end_vn1070);
V1071:VNPU6_6 port map (start_vn,clk,rst,Lc1071,C99V1071,C207V1071,C512V1071,C828V1071,C903V1071,C1141V1071,V1071C99,V1071C207,V1071C512,V1071C828,V1071C903,V1071C1141,SI1071,end_vn1071);
V1072:VNPU6_6 port map (start_vn,clk,rst,Lc1072,C100V1072,C208V1072,C513V1072,C829V1072,C904V1072,C1142V1072,V1072C100,V1072C208,V1072C513,V1072C829,V1072C904,V1072C1142,SI1072,end_vn1072);
V1073:VNPU6_6 port map (start_vn,clk,rst,Lc1073,C101V1073,C209V1073,C514V1073,C830V1073,C905V1073,C1143V1073,V1073C101,V1073C209,V1073C514,V1073C830,V1073C905,V1073C1143,SI1073,end_vn1073);
V1074:VNPU6_6 port map (start_vn,clk,rst,Lc1074,C102V1074,C210V1074,C515V1074,C831V1074,C906V1074,C1144V1074,V1074C102,V1074C210,V1074C515,V1074C831,V1074C906,V1074C1144,SI1074,end_vn1074);
V1075:VNPU6_6 port map (start_vn,clk,rst,Lc1075,C103V1075,C211V1075,C516V1075,C832V1075,C907V1075,C1145V1075,V1075C103,V1075C211,V1075C516,V1075C832,V1075C907,V1075C1145,SI1075,end_vn1075);
V1076:VNPU6_6 port map (start_vn,clk,rst,Lc1076,C104V1076,C212V1076,C517V1076,C833V1076,C908V1076,C1146V1076,V1076C104,V1076C212,V1076C517,V1076C833,V1076C908,V1076C1146,SI1076,end_vn1076);
V1077:VNPU6_6 port map (start_vn,clk,rst,Lc1077,C105V1077,C213V1077,C518V1077,C834V1077,C909V1077,C1147V1077,V1077C105,V1077C213,V1077C518,V1077C834,V1077C909,V1077C1147,SI1077,end_vn1077);
V1078:VNPU6_6 port map (start_vn,clk,rst,Lc1078,C106V1078,C214V1078,C519V1078,C835V1078,C910V1078,C1148V1078,V1078C106,V1078C214,V1078C519,V1078C835,V1078C910,V1078C1148,SI1078,end_vn1078);
V1079:VNPU6_6 port map (start_vn,clk,rst,Lc1079,C107V1079,C215V1079,C520V1079,C836V1079,C911V1079,C1149V1079,V1079C107,V1079C215,V1079C520,V1079C836,V1079C911,V1079C1149,SI1079,end_vn1079);
V1080:VNPU6_6 port map (start_vn,clk,rst,Lc1080,C108V1080,C216V1080,C521V1080,C837V1080,C912V1080,C1150V1080,V1080C108,V1080C216,V1080C521,V1080C837,V1080C912,V1080C1150,SI1080,end_vn1080);
V1081:VNPU6_6 port map (start_vn,clk,rst,Lc1081,C109V1081,C217V1081,C522V1081,C838V1081,C913V1081,C1151V1081,V1081C109,V1081C217,V1081C522,V1081C838,V1081C913,V1081C1151,SI1081,end_vn1081);
V1082:VNPU6_6 port map (start_vn,clk,rst,Lc1082,C110V1082,C218V1082,C523V1082,C839V1082,C914V1082,C1152V1082,V1082C110,V1082C218,V1082C523,V1082C839,V1082C914,V1082C1152,SI1082,end_vn1082);
V1083:VNPU6_6 port map (start_vn,clk,rst,Lc1083,C111V1083,C219V1083,C524V1083,C840V1083,C915V1083,C1057V1083,V1083C111,V1083C219,V1083C524,V1083C840,V1083C915,V1083C1057,SI1083,end_vn1083);
V1084:VNPU6_6 port map (start_vn,clk,rst,Lc1084,C112V1084,C220V1084,C525V1084,C841V1084,C916V1084,C1058V1084,V1084C112,V1084C220,V1084C525,V1084C841,V1084C916,V1084C1058,SI1084,end_vn1084);
V1085:VNPU6_6 port map (start_vn,clk,rst,Lc1085,C113V1085,C221V1085,C526V1085,C842V1085,C917V1085,C1059V1085,V1085C113,V1085C221,V1085C526,V1085C842,V1085C917,V1085C1059,SI1085,end_vn1085);
V1086:VNPU6_6 port map (start_vn,clk,rst,Lc1086,C114V1086,C222V1086,C527V1086,C843V1086,C918V1086,C1060V1086,V1086C114,V1086C222,V1086C527,V1086C843,V1086C918,V1086C1060,SI1086,end_vn1086);
V1087:VNPU6_6 port map (start_vn,clk,rst,Lc1087,C115V1087,C223V1087,C528V1087,C844V1087,C919V1087,C1061V1087,V1087C115,V1087C223,V1087C528,V1087C844,V1087C919,V1087C1061,SI1087,end_vn1087);
V1088:VNPU6_6 port map (start_vn,clk,rst,Lc1088,C116V1088,C224V1088,C529V1088,C845V1088,C920V1088,C1062V1088,V1088C116,V1088C224,V1088C529,V1088C845,V1088C920,V1088C1062,SI1088,end_vn1088);
V1089:VNPU6_6 port map (start_vn,clk,rst,Lc1089,C117V1089,C225V1089,C530V1089,C846V1089,C921V1089,C1063V1089,V1089C117,V1089C225,V1089C530,V1089C846,V1089C921,V1089C1063,SI1089,end_vn1089);
V1090:VNPU6_6 port map (start_vn,clk,rst,Lc1090,C118V1090,C226V1090,C531V1090,C847V1090,C922V1090,C1064V1090,V1090C118,V1090C226,V1090C531,V1090C847,V1090C922,V1090C1064,SI1090,end_vn1090);
V1091:VNPU6_6 port map (start_vn,clk,rst,Lc1091,C119V1091,C227V1091,C532V1091,C848V1091,C923V1091,C1065V1091,V1091C119,V1091C227,V1091C532,V1091C848,V1091C923,V1091C1065,SI1091,end_vn1091);
V1092:VNPU6_6 port map (start_vn,clk,rst,Lc1092,C120V1092,C228V1092,C533V1092,C849V1092,C924V1092,C1066V1092,V1092C120,V1092C228,V1092C533,V1092C849,V1092C924,V1092C1066,SI1092,end_vn1092);
V1093:VNPU6_6 port map (start_vn,clk,rst,Lc1093,C121V1093,C229V1093,C534V1093,C850V1093,C925V1093,C1067V1093,V1093C121,V1093C229,V1093C534,V1093C850,V1093C925,V1093C1067,SI1093,end_vn1093);
V1094:VNPU6_6 port map (start_vn,clk,rst,Lc1094,C122V1094,C230V1094,C535V1094,C851V1094,C926V1094,C1068V1094,V1094C122,V1094C230,V1094C535,V1094C851,V1094C926,V1094C1068,SI1094,end_vn1094);
V1095:VNPU6_6 port map (start_vn,clk,rst,Lc1095,C123V1095,C231V1095,C536V1095,C852V1095,C927V1095,C1069V1095,V1095C123,V1095C231,V1095C536,V1095C852,V1095C927,V1095C1069,SI1095,end_vn1095);
V1096:VNPU6_6 port map (start_vn,clk,rst,Lc1096,C124V1096,C232V1096,C537V1096,C853V1096,C928V1096,C1070V1096,V1096C124,V1096C232,V1096C537,V1096C853,V1096C928,V1096C1070,SI1096,end_vn1096);
V1097:VNPU6_6 port map (start_vn,clk,rst,Lc1097,C125V1097,C233V1097,C538V1097,C854V1097,C929V1097,C1071V1097,V1097C125,V1097C233,V1097C538,V1097C854,V1097C929,V1097C1071,SI1097,end_vn1097);
V1098:VNPU6_6 port map (start_vn,clk,rst,Lc1098,C126V1098,C234V1098,C539V1098,C855V1098,C930V1098,C1072V1098,V1098C126,V1098C234,V1098C539,V1098C855,V1098C930,V1098C1072,SI1098,end_vn1098);
V1099:VNPU6_6 port map (start_vn,clk,rst,Lc1099,C127V1099,C235V1099,C540V1099,C856V1099,C931V1099,C1073V1099,V1099C127,V1099C235,V1099C540,V1099C856,V1099C931,V1099C1073,SI1099,end_vn1099);
V1100:VNPU6_6 port map (start_vn,clk,rst,Lc1100,C128V1100,C236V1100,C541V1100,C857V1100,C932V1100,C1074V1100,V1100C128,V1100C236,V1100C541,V1100C857,V1100C932,V1100C1074,SI1100,end_vn1100);
V1101:VNPU6_6 port map (start_vn,clk,rst,Lc1101,C129V1101,C237V1101,C542V1101,C858V1101,C933V1101,C1075V1101,V1101C129,V1101C237,V1101C542,V1101C858,V1101C933,V1101C1075,SI1101,end_vn1101);
V1102:VNPU6_6 port map (start_vn,clk,rst,Lc1102,C130V1102,C238V1102,C543V1102,C859V1102,C934V1102,C1076V1102,V1102C130,V1102C238,V1102C543,V1102C859,V1102C934,V1102C1076,SI1102,end_vn1102);
V1103:VNPU6_6 port map (start_vn,clk,rst,Lc1103,C131V1103,C239V1103,C544V1103,C860V1103,C935V1103,C1077V1103,V1103C131,V1103C239,V1103C544,V1103C860,V1103C935,V1103C1077,SI1103,end_vn1103);
V1104:VNPU6_6 port map (start_vn,clk,rst,Lc1104,C132V1104,C240V1104,C545V1104,C861V1104,C936V1104,C1078V1104,V1104C132,V1104C240,V1104C545,V1104C861,V1104C936,V1104C1078,SI1104,end_vn1104);
V1105:VNPU6_6 port map (start_vn,clk,rst,Lc1105,C133V1105,C241V1105,C546V1105,C862V1105,C937V1105,C1079V1105,V1105C133,V1105C241,V1105C546,V1105C862,V1105C937,V1105C1079,SI1105,end_vn1105);
V1106:VNPU6_6 port map (start_vn,clk,rst,Lc1106,C134V1106,C242V1106,C547V1106,C863V1106,C938V1106,C1080V1106,V1106C134,V1106C242,V1106C547,V1106C863,V1106C938,V1106C1080,SI1106,end_vn1106);
V1107:VNPU6_6 port map (start_vn,clk,rst,Lc1107,C135V1107,C243V1107,C548V1107,C864V1107,C939V1107,C1081V1107,V1107C135,V1107C243,V1107C548,V1107C864,V1107C939,V1107C1081,SI1107,end_vn1107);
V1108:VNPU6_6 port map (start_vn,clk,rst,Lc1108,C136V1108,C244V1108,C549V1108,C769V1108,C940V1108,C1082V1108,V1108C136,V1108C244,V1108C549,V1108C769,V1108C940,V1108C1082,SI1108,end_vn1108);
V1109:VNPU6_6 port map (start_vn,clk,rst,Lc1109,C137V1109,C245V1109,C550V1109,C770V1109,C941V1109,C1083V1109,V1109C137,V1109C245,V1109C550,V1109C770,V1109C941,V1109C1083,SI1109,end_vn1109);
V1110:VNPU6_6 port map (start_vn,clk,rst,Lc1110,C138V1110,C246V1110,C551V1110,C771V1110,C942V1110,C1084V1110,V1110C138,V1110C246,V1110C551,V1110C771,V1110C942,V1110C1084,SI1110,end_vn1110);
V1111:VNPU6_6 port map (start_vn,clk,rst,Lc1111,C139V1111,C247V1111,C552V1111,C772V1111,C943V1111,C1085V1111,V1111C139,V1111C247,V1111C552,V1111C772,V1111C943,V1111C1085,SI1111,end_vn1111);
V1112:VNPU6_6 port map (start_vn,clk,rst,Lc1112,C140V1112,C248V1112,C553V1112,C773V1112,C944V1112,C1086V1112,V1112C140,V1112C248,V1112C553,V1112C773,V1112C944,V1112C1086,SI1112,end_vn1112);
V1113:VNPU6_6 port map (start_vn,clk,rst,Lc1113,C141V1113,C249V1113,C554V1113,C774V1113,C945V1113,C1087V1113,V1113C141,V1113C249,V1113C554,V1113C774,V1113C945,V1113C1087,SI1113,end_vn1113);
V1114:VNPU6_6 port map (start_vn,clk,rst,Lc1114,C142V1114,C250V1114,C555V1114,C775V1114,C946V1114,C1088V1114,V1114C142,V1114C250,V1114C555,V1114C775,V1114C946,V1114C1088,SI1114,end_vn1114);
V1115:VNPU6_6 port map (start_vn,clk,rst,Lc1115,C143V1115,C251V1115,C556V1115,C776V1115,C947V1115,C1089V1115,V1115C143,V1115C251,V1115C556,V1115C776,V1115C947,V1115C1089,SI1115,end_vn1115);
V1116:VNPU6_6 port map (start_vn,clk,rst,Lc1116,C144V1116,C252V1116,C557V1116,C777V1116,C948V1116,C1090V1116,V1116C144,V1116C252,V1116C557,V1116C777,V1116C948,V1116C1090,SI1116,end_vn1116);
V1117:VNPU6_6 port map (start_vn,clk,rst,Lc1117,C145V1117,C253V1117,C558V1117,C778V1117,C949V1117,C1091V1117,V1117C145,V1117C253,V1117C558,V1117C778,V1117C949,V1117C1091,SI1117,end_vn1117);
V1118:VNPU6_6 port map (start_vn,clk,rst,Lc1118,C146V1118,C254V1118,C559V1118,C779V1118,C950V1118,C1092V1118,V1118C146,V1118C254,V1118C559,V1118C779,V1118C950,V1118C1092,SI1118,end_vn1118);
V1119:VNPU6_6 port map (start_vn,clk,rst,Lc1119,C147V1119,C255V1119,C560V1119,C780V1119,C951V1119,C1093V1119,V1119C147,V1119C255,V1119C560,V1119C780,V1119C951,V1119C1093,SI1119,end_vn1119);
V1120:VNPU6_6 port map (start_vn,clk,rst,Lc1120,C148V1120,C256V1120,C561V1120,C781V1120,C952V1120,C1094V1120,V1120C148,V1120C256,V1120C561,V1120C781,V1120C952,V1120C1094,SI1120,end_vn1120);
V1121:VNPU6_6 port map (start_vn,clk,rst,Lc1121,C149V1121,C257V1121,C562V1121,C782V1121,C953V1121,C1095V1121,V1121C149,V1121C257,V1121C562,V1121C782,V1121C953,V1121C1095,SI1121,end_vn1121);
V1122:VNPU6_6 port map (start_vn,clk,rst,Lc1122,C150V1122,C258V1122,C563V1122,C783V1122,C954V1122,C1096V1122,V1122C150,V1122C258,V1122C563,V1122C783,V1122C954,V1122C1096,SI1122,end_vn1122);
V1123:VNPU6_6 port map (start_vn,clk,rst,Lc1123,C151V1123,C259V1123,C564V1123,C784V1123,C955V1123,C1097V1123,V1123C151,V1123C259,V1123C564,V1123C784,V1123C955,V1123C1097,SI1123,end_vn1123);
V1124:VNPU6_6 port map (start_vn,clk,rst,Lc1124,C152V1124,C260V1124,C565V1124,C785V1124,C956V1124,C1098V1124,V1124C152,V1124C260,V1124C565,V1124C785,V1124C956,V1124C1098,SI1124,end_vn1124);
V1125:VNPU6_6 port map (start_vn,clk,rst,Lc1125,C153V1125,C261V1125,C566V1125,C786V1125,C957V1125,C1099V1125,V1125C153,V1125C261,V1125C566,V1125C786,V1125C957,V1125C1099,SI1125,end_vn1125);
V1126:VNPU6_6 port map (start_vn,clk,rst,Lc1126,C154V1126,C262V1126,C567V1126,C787V1126,C958V1126,C1100V1126,V1126C154,V1126C262,V1126C567,V1126C787,V1126C958,V1126C1100,SI1126,end_vn1126);
V1127:VNPU6_6 port map (start_vn,clk,rst,Lc1127,C155V1127,C263V1127,C568V1127,C788V1127,C959V1127,C1101V1127,V1127C155,V1127C263,V1127C568,V1127C788,V1127C959,V1127C1101,SI1127,end_vn1127);
V1128:VNPU6_6 port map (start_vn,clk,rst,Lc1128,C156V1128,C264V1128,C569V1128,C789V1128,C960V1128,C1102V1128,V1128C156,V1128C264,V1128C569,V1128C789,V1128C960,V1128C1102,SI1128,end_vn1128);
V1129:VNPU6_6 port map (start_vn,clk,rst,Lc1129,C157V1129,C265V1129,C570V1129,C790V1129,C865V1129,C1103V1129,V1129C157,V1129C265,V1129C570,V1129C790,V1129C865,V1129C1103,SI1129,end_vn1129);
V1130:VNPU6_6 port map (start_vn,clk,rst,Lc1130,C158V1130,C266V1130,C571V1130,C791V1130,C866V1130,C1104V1130,V1130C158,V1130C266,V1130C571,V1130C791,V1130C866,V1130C1104,SI1130,end_vn1130);
V1131:VNPU6_6 port map (start_vn,clk,rst,Lc1131,C159V1131,C267V1131,C572V1131,C792V1131,C867V1131,C1105V1131,V1131C159,V1131C267,V1131C572,V1131C792,V1131C867,V1131C1105,SI1131,end_vn1131);
V1132:VNPU6_6 port map (start_vn,clk,rst,Lc1132,C160V1132,C268V1132,C573V1132,C793V1132,C868V1132,C1106V1132,V1132C160,V1132C268,V1132C573,V1132C793,V1132C868,V1132C1106,SI1132,end_vn1132);
V1133:VNPU6_6 port map (start_vn,clk,rst,Lc1133,C161V1133,C269V1133,C574V1133,C794V1133,C869V1133,C1107V1133,V1133C161,V1133C269,V1133C574,V1133C794,V1133C869,V1133C1107,SI1133,end_vn1133);
V1134:VNPU6_6 port map (start_vn,clk,rst,Lc1134,C162V1134,C270V1134,C575V1134,C795V1134,C870V1134,C1108V1134,V1134C162,V1134C270,V1134C575,V1134C795,V1134C870,V1134C1108,SI1134,end_vn1134);
V1135:VNPU6_6 port map (start_vn,clk,rst,Lc1135,C163V1135,C271V1135,C576V1135,C796V1135,C871V1135,C1109V1135,V1135C163,V1135C271,V1135C576,V1135C796,V1135C871,V1135C1109,SI1135,end_vn1135);
V1136:VNPU6_6 port map (start_vn,clk,rst,Lc1136,C164V1136,C272V1136,C481V1136,C797V1136,C872V1136,C1110V1136,V1136C164,V1136C272,V1136C481,V1136C797,V1136C872,V1136C1110,SI1136,end_vn1136);
V1137:VNPU6_6 port map (start_vn,clk,rst,Lc1137,C165V1137,C273V1137,C482V1137,C798V1137,C873V1137,C1111V1137,V1137C165,V1137C273,V1137C482,V1137C798,V1137C873,V1137C1111,SI1137,end_vn1137);
V1138:VNPU6_6 port map (start_vn,clk,rst,Lc1138,C166V1138,C274V1138,C483V1138,C799V1138,C874V1138,C1112V1138,V1138C166,V1138C274,V1138C483,V1138C799,V1138C874,V1138C1112,SI1138,end_vn1138);
V1139:VNPU6_6 port map (start_vn,clk,rst,Lc1139,C167V1139,C275V1139,C484V1139,C800V1139,C875V1139,C1113V1139,V1139C167,V1139C275,V1139C484,V1139C800,V1139C875,V1139C1113,SI1139,end_vn1139);
V1140:VNPU6_6 port map (start_vn,clk,rst,Lc1140,C168V1140,C276V1140,C485V1140,C801V1140,C876V1140,C1114V1140,V1140C168,V1140C276,V1140C485,V1140C801,V1140C876,V1140C1114,SI1140,end_vn1140);
V1141:VNPU6_6 port map (start_vn,clk,rst,Lc1141,C169V1141,C277V1141,C486V1141,C802V1141,C877V1141,C1115V1141,V1141C169,V1141C277,V1141C486,V1141C802,V1141C877,V1141C1115,SI1141,end_vn1141);
V1142:VNPU6_6 port map (start_vn,clk,rst,Lc1142,C170V1142,C278V1142,C487V1142,C803V1142,C878V1142,C1116V1142,V1142C170,V1142C278,V1142C487,V1142C803,V1142C878,V1142C1116,SI1142,end_vn1142);
V1143:VNPU6_6 port map (start_vn,clk,rst,Lc1143,C171V1143,C279V1143,C488V1143,C804V1143,C879V1143,C1117V1143,V1143C171,V1143C279,V1143C488,V1143C804,V1143C879,V1143C1117,SI1143,end_vn1143);
V1144:VNPU6_6 port map (start_vn,clk,rst,Lc1144,C172V1144,C280V1144,C489V1144,C805V1144,C880V1144,C1118V1144,V1144C172,V1144C280,V1144C489,V1144C805,V1144C880,V1144C1118,SI1144,end_vn1144);
V1145:VNPU6_6 port map (start_vn,clk,rst,Lc1145,C173V1145,C281V1145,C490V1145,C806V1145,C881V1145,C1119V1145,V1145C173,V1145C281,V1145C490,V1145C806,V1145C881,V1145C1119,SI1145,end_vn1145);
V1146:VNPU6_6 port map (start_vn,clk,rst,Lc1146,C174V1146,C282V1146,C491V1146,C807V1146,C882V1146,C1120V1146,V1146C174,V1146C282,V1146C491,V1146C807,V1146C882,V1146C1120,SI1146,end_vn1146);
V1147:VNPU6_6 port map (start_vn,clk,rst,Lc1147,C175V1147,C283V1147,C492V1147,C808V1147,C883V1147,C1121V1147,V1147C175,V1147C283,V1147C492,V1147C808,V1147C883,V1147C1121,SI1147,end_vn1147);
V1148:VNPU6_6 port map (start_vn,clk,rst,Lc1148,C176V1148,C284V1148,C493V1148,C809V1148,C884V1148,C1122V1148,V1148C176,V1148C284,V1148C493,V1148C809,V1148C884,V1148C1122,SI1148,end_vn1148);
V1149:VNPU6_6 port map (start_vn,clk,rst,Lc1149,C177V1149,C285V1149,C494V1149,C810V1149,C885V1149,C1123V1149,V1149C177,V1149C285,V1149C494,V1149C810,V1149C885,V1149C1123,SI1149,end_vn1149);
V1150:VNPU6_6 port map (start_vn,clk,rst,Lc1150,C178V1150,C286V1150,C495V1150,C811V1150,C886V1150,C1124V1150,V1150C178,V1150C286,V1150C495,V1150C811,V1150C886,V1150C1124,SI1150,end_vn1150);
V1151:VNPU6_6 port map (start_vn,clk,rst,Lc1151,C179V1151,C287V1151,C496V1151,C812V1151,C887V1151,C1125V1151,V1151C179,V1151C287,V1151C496,V1151C812,V1151C887,V1151C1125,SI1151,end_vn1151);
V1152:VNPU6_6 port map (start_vn,clk,rst,Lc1152,C180V1152,C288V1152,C497V1152,C813V1152,C888V1152,C1126V1152,V1152C180,V1152C288,V1152C497,V1152C813,V1152C888,V1152C1126,SI1152,end_vn1152);
V1153:VNPU3_3 port map (start_vn,clk,rst,Lc1153,C90V1153,C481V1153,C1146V1153,V1153C90,V1153C481,V1153C1146,SI1153,end_vn1153);
V1154:VNPU3_3 port map (start_vn,clk,rst,Lc1154,C91V1154,C482V1154,C1147V1154,V1154C91,V1154C482,V1154C1147,SI1154,end_vn1154);
V1155:VNPU3_3 port map (start_vn,clk,rst,Lc1155,C92V1155,C483V1155,C1148V1155,V1155C92,V1155C483,V1155C1148,SI1155,end_vn1155);
V1156:VNPU3_3 port map (start_vn,clk,rst,Lc1156,C93V1156,C484V1156,C1149V1156,V1156C93,V1156C484,V1156C1149,SI1156,end_vn1156);
V1157:VNPU3_3 port map (start_vn,clk,rst,Lc1157,C94V1157,C485V1157,C1150V1157,V1157C94,V1157C485,V1157C1150,SI1157,end_vn1157);
V1158:VNPU3_3 port map (start_vn,clk,rst,Lc1158,C95V1158,C486V1158,C1151V1158,V1158C95,V1158C486,V1158C1151,SI1158,end_vn1158);
V1159:VNPU3_3 port map (start_vn,clk,rst,Lc1159,C96V1159,C487V1159,C1152V1159,V1159C96,V1159C487,V1159C1152,SI1159,end_vn1159);
V1160:VNPU3_3 port map (start_vn,clk,rst,Lc1160,C1V1160,C488V1160,C1057V1160,V1160C1,V1160C488,V1160C1057,SI1160,end_vn1160);
V1161:VNPU3_3 port map (start_vn,clk,rst,Lc1161,C2V1161,C489V1161,C1058V1161,V1161C2,V1161C489,V1161C1058,SI1161,end_vn1161);
V1162:VNPU3_3 port map (start_vn,clk,rst,Lc1162,C3V1162,C490V1162,C1059V1162,V1162C3,V1162C490,V1162C1059,SI1162,end_vn1162);
V1163:VNPU3_3 port map (start_vn,clk,rst,Lc1163,C4V1163,C491V1163,C1060V1163,V1163C4,V1163C491,V1163C1060,SI1163,end_vn1163);
V1164:VNPU3_3 port map (start_vn,clk,rst,Lc1164,C5V1164,C492V1164,C1061V1164,V1164C5,V1164C492,V1164C1061,SI1164,end_vn1164);
V1165:VNPU3_3 port map (start_vn,clk,rst,Lc1165,C6V1165,C493V1165,C1062V1165,V1165C6,V1165C493,V1165C1062,SI1165,end_vn1165);
V1166:VNPU3_3 port map (start_vn,clk,rst,Lc1166,C7V1166,C494V1166,C1063V1166,V1166C7,V1166C494,V1166C1063,SI1166,end_vn1166);
V1167:VNPU3_3 port map (start_vn,clk,rst,Lc1167,C8V1167,C495V1167,C1064V1167,V1167C8,V1167C495,V1167C1064,SI1167,end_vn1167);
V1168:VNPU3_3 port map (start_vn,clk,rst,Lc1168,C9V1168,C496V1168,C1065V1168,V1168C9,V1168C496,V1168C1065,SI1168,end_vn1168);
V1169:VNPU3_3 port map (start_vn,clk,rst,Lc1169,C10V1169,C497V1169,C1066V1169,V1169C10,V1169C497,V1169C1066,SI1169,end_vn1169);
V1170:VNPU3_3 port map (start_vn,clk,rst,Lc1170,C11V1170,C498V1170,C1067V1170,V1170C11,V1170C498,V1170C1067,SI1170,end_vn1170);
V1171:VNPU3_3 port map (start_vn,clk,rst,Lc1171,C12V1171,C499V1171,C1068V1171,V1171C12,V1171C499,V1171C1068,SI1171,end_vn1171);
V1172:VNPU3_3 port map (start_vn,clk,rst,Lc1172,C13V1172,C500V1172,C1069V1172,V1172C13,V1172C500,V1172C1069,SI1172,end_vn1172);
V1173:VNPU3_3 port map (start_vn,clk,rst,Lc1173,C14V1173,C501V1173,C1070V1173,V1173C14,V1173C501,V1173C1070,SI1173,end_vn1173);
V1174:VNPU3_3 port map (start_vn,clk,rst,Lc1174,C15V1174,C502V1174,C1071V1174,V1174C15,V1174C502,V1174C1071,SI1174,end_vn1174);
V1175:VNPU3_3 port map (start_vn,clk,rst,Lc1175,C16V1175,C503V1175,C1072V1175,V1175C16,V1175C503,V1175C1072,SI1175,end_vn1175);
V1176:VNPU3_3 port map (start_vn,clk,rst,Lc1176,C17V1176,C504V1176,C1073V1176,V1176C17,V1176C504,V1176C1073,SI1176,end_vn1176);
V1177:VNPU3_3 port map (start_vn,clk,rst,Lc1177,C18V1177,C505V1177,C1074V1177,V1177C18,V1177C505,V1177C1074,SI1177,end_vn1177);
V1178:VNPU3_3 port map (start_vn,clk,rst,Lc1178,C19V1178,C506V1178,C1075V1178,V1178C19,V1178C506,V1178C1075,SI1178,end_vn1178);
V1179:VNPU3_3 port map (start_vn,clk,rst,Lc1179,C20V1179,C507V1179,C1076V1179,V1179C20,V1179C507,V1179C1076,SI1179,end_vn1179);
V1180:VNPU3_3 port map (start_vn,clk,rst,Lc1180,C21V1180,C508V1180,C1077V1180,V1180C21,V1180C508,V1180C1077,SI1180,end_vn1180);
V1181:VNPU3_3 port map (start_vn,clk,rst,Lc1181,C22V1181,C509V1181,C1078V1181,V1181C22,V1181C509,V1181C1078,SI1181,end_vn1181);
V1182:VNPU3_3 port map (start_vn,clk,rst,Lc1182,C23V1182,C510V1182,C1079V1182,V1182C23,V1182C510,V1182C1079,SI1182,end_vn1182);
V1183:VNPU3_3 port map (start_vn,clk,rst,Lc1183,C24V1183,C511V1183,C1080V1183,V1183C24,V1183C511,V1183C1080,SI1183,end_vn1183);
V1184:VNPU3_3 port map (start_vn,clk,rst,Lc1184,C25V1184,C512V1184,C1081V1184,V1184C25,V1184C512,V1184C1081,SI1184,end_vn1184);
V1185:VNPU3_3 port map (start_vn,clk,rst,Lc1185,C26V1185,C513V1185,C1082V1185,V1185C26,V1185C513,V1185C1082,SI1185,end_vn1185);
V1186:VNPU3_3 port map (start_vn,clk,rst,Lc1186,C27V1186,C514V1186,C1083V1186,V1186C27,V1186C514,V1186C1083,SI1186,end_vn1186);
V1187:VNPU3_3 port map (start_vn,clk,rst,Lc1187,C28V1187,C515V1187,C1084V1187,V1187C28,V1187C515,V1187C1084,SI1187,end_vn1187);
V1188:VNPU3_3 port map (start_vn,clk,rst,Lc1188,C29V1188,C516V1188,C1085V1188,V1188C29,V1188C516,V1188C1085,SI1188,end_vn1188);
V1189:VNPU3_3 port map (start_vn,clk,rst,Lc1189,C30V1189,C517V1189,C1086V1189,V1189C30,V1189C517,V1189C1086,SI1189,end_vn1189);
V1190:VNPU3_3 port map (start_vn,clk,rst,Lc1190,C31V1190,C518V1190,C1087V1190,V1190C31,V1190C518,V1190C1087,SI1190,end_vn1190);
V1191:VNPU3_3 port map (start_vn,clk,rst,Lc1191,C32V1191,C519V1191,C1088V1191,V1191C32,V1191C519,V1191C1088,SI1191,end_vn1191);
V1192:VNPU3_3 port map (start_vn,clk,rst,Lc1192,C33V1192,C520V1192,C1089V1192,V1192C33,V1192C520,V1192C1089,SI1192,end_vn1192);
V1193:VNPU3_3 port map (start_vn,clk,rst,Lc1193,C34V1193,C521V1193,C1090V1193,V1193C34,V1193C521,V1193C1090,SI1193,end_vn1193);
V1194:VNPU3_3 port map (start_vn,clk,rst,Lc1194,C35V1194,C522V1194,C1091V1194,V1194C35,V1194C522,V1194C1091,SI1194,end_vn1194);
V1195:VNPU3_3 port map (start_vn,clk,rst,Lc1195,C36V1195,C523V1195,C1092V1195,V1195C36,V1195C523,V1195C1092,SI1195,end_vn1195);
V1196:VNPU3_3 port map (start_vn,clk,rst,Lc1196,C37V1196,C524V1196,C1093V1196,V1196C37,V1196C524,V1196C1093,SI1196,end_vn1196);
V1197:VNPU3_3 port map (start_vn,clk,rst,Lc1197,C38V1197,C525V1197,C1094V1197,V1197C38,V1197C525,V1197C1094,SI1197,end_vn1197);
V1198:VNPU3_3 port map (start_vn,clk,rst,Lc1198,C39V1198,C526V1198,C1095V1198,V1198C39,V1198C526,V1198C1095,SI1198,end_vn1198);
V1199:VNPU3_3 port map (start_vn,clk,rst,Lc1199,C40V1199,C527V1199,C1096V1199,V1199C40,V1199C527,V1199C1096,SI1199,end_vn1199);
V1200:VNPU3_3 port map (start_vn,clk,rst,Lc1200,C41V1200,C528V1200,C1097V1200,V1200C41,V1200C528,V1200C1097,SI1200,end_vn1200);
V1201:VNPU3_3 port map (start_vn,clk,rst,Lc1201,C42V1201,C529V1201,C1098V1201,V1201C42,V1201C529,V1201C1098,SI1201,end_vn1201);
V1202:VNPU3_3 port map (start_vn,clk,rst,Lc1202,C43V1202,C530V1202,C1099V1202,V1202C43,V1202C530,V1202C1099,SI1202,end_vn1202);
V1203:VNPU3_3 port map (start_vn,clk,rst,Lc1203,C44V1203,C531V1203,C1100V1203,V1203C44,V1203C531,V1203C1100,SI1203,end_vn1203);
V1204:VNPU3_3 port map (start_vn,clk,rst,Lc1204,C45V1204,C532V1204,C1101V1204,V1204C45,V1204C532,V1204C1101,SI1204,end_vn1204);
V1205:VNPU3_3 port map (start_vn,clk,rst,Lc1205,C46V1205,C533V1205,C1102V1205,V1205C46,V1205C533,V1205C1102,SI1205,end_vn1205);
V1206:VNPU3_3 port map (start_vn,clk,rst,Lc1206,C47V1206,C534V1206,C1103V1206,V1206C47,V1206C534,V1206C1103,SI1206,end_vn1206);
V1207:VNPU3_3 port map (start_vn,clk,rst,Lc1207,C48V1207,C535V1207,C1104V1207,V1207C48,V1207C535,V1207C1104,SI1207,end_vn1207);
V1208:VNPU3_3 port map (start_vn,clk,rst,Lc1208,C49V1208,C536V1208,C1105V1208,V1208C49,V1208C536,V1208C1105,SI1208,end_vn1208);
V1209:VNPU3_3 port map (start_vn,clk,rst,Lc1209,C50V1209,C537V1209,C1106V1209,V1209C50,V1209C537,V1209C1106,SI1209,end_vn1209);
V1210:VNPU3_3 port map (start_vn,clk,rst,Lc1210,C51V1210,C538V1210,C1107V1210,V1210C51,V1210C538,V1210C1107,SI1210,end_vn1210);
V1211:VNPU3_3 port map (start_vn,clk,rst,Lc1211,C52V1211,C539V1211,C1108V1211,V1211C52,V1211C539,V1211C1108,SI1211,end_vn1211);
V1212:VNPU3_3 port map (start_vn,clk,rst,Lc1212,C53V1212,C540V1212,C1109V1212,V1212C53,V1212C540,V1212C1109,SI1212,end_vn1212);
V1213:VNPU3_3 port map (start_vn,clk,rst,Lc1213,C54V1213,C541V1213,C1110V1213,V1213C54,V1213C541,V1213C1110,SI1213,end_vn1213);
V1214:VNPU3_3 port map (start_vn,clk,rst,Lc1214,C55V1214,C542V1214,C1111V1214,V1214C55,V1214C542,V1214C1111,SI1214,end_vn1214);
V1215:VNPU3_3 port map (start_vn,clk,rst,Lc1215,C56V1215,C543V1215,C1112V1215,V1215C56,V1215C543,V1215C1112,SI1215,end_vn1215);
V1216:VNPU3_3 port map (start_vn,clk,rst,Lc1216,C57V1216,C544V1216,C1113V1216,V1216C57,V1216C544,V1216C1113,SI1216,end_vn1216);
V1217:VNPU3_3 port map (start_vn,clk,rst,Lc1217,C58V1217,C545V1217,C1114V1217,V1217C58,V1217C545,V1217C1114,SI1217,end_vn1217);
V1218:VNPU3_3 port map (start_vn,clk,rst,Lc1218,C59V1218,C546V1218,C1115V1218,V1218C59,V1218C546,V1218C1115,SI1218,end_vn1218);
V1219:VNPU3_3 port map (start_vn,clk,rst,Lc1219,C60V1219,C547V1219,C1116V1219,V1219C60,V1219C547,V1219C1116,SI1219,end_vn1219);
V1220:VNPU3_3 port map (start_vn,clk,rst,Lc1220,C61V1220,C548V1220,C1117V1220,V1220C61,V1220C548,V1220C1117,SI1220,end_vn1220);
V1221:VNPU3_3 port map (start_vn,clk,rst,Lc1221,C62V1221,C549V1221,C1118V1221,V1221C62,V1221C549,V1221C1118,SI1221,end_vn1221);
V1222:VNPU3_3 port map (start_vn,clk,rst,Lc1222,C63V1222,C550V1222,C1119V1222,V1222C63,V1222C550,V1222C1119,SI1222,end_vn1222);
V1223:VNPU3_3 port map (start_vn,clk,rst,Lc1223,C64V1223,C551V1223,C1120V1223,V1223C64,V1223C551,V1223C1120,SI1223,end_vn1223);
V1224:VNPU3_3 port map (start_vn,clk,rst,Lc1224,C65V1224,C552V1224,C1121V1224,V1224C65,V1224C552,V1224C1121,SI1224,end_vn1224);
V1225:VNPU3_3 port map (start_vn,clk,rst,Lc1225,C66V1225,C553V1225,C1122V1225,V1225C66,V1225C553,V1225C1122,SI1225,end_vn1225);
V1226:VNPU3_3 port map (start_vn,clk,rst,Lc1226,C67V1226,C554V1226,C1123V1226,V1226C67,V1226C554,V1226C1123,SI1226,end_vn1226);
V1227:VNPU3_3 port map (start_vn,clk,rst,Lc1227,C68V1227,C555V1227,C1124V1227,V1227C68,V1227C555,V1227C1124,SI1227,end_vn1227);
V1228:VNPU3_3 port map (start_vn,clk,rst,Lc1228,C69V1228,C556V1228,C1125V1228,V1228C69,V1228C556,V1228C1125,SI1228,end_vn1228);
V1229:VNPU3_3 port map (start_vn,clk,rst,Lc1229,C70V1229,C557V1229,C1126V1229,V1229C70,V1229C557,V1229C1126,SI1229,end_vn1229);
V1230:VNPU3_3 port map (start_vn,clk,rst,Lc1230,C71V1230,C558V1230,C1127V1230,V1230C71,V1230C558,V1230C1127,SI1230,end_vn1230);
V1231:VNPU3_3 port map (start_vn,clk,rst,Lc1231,C72V1231,C559V1231,C1128V1231,V1231C72,V1231C559,V1231C1128,SI1231,end_vn1231);
V1232:VNPU3_3 port map (start_vn,clk,rst,Lc1232,C73V1232,C560V1232,C1129V1232,V1232C73,V1232C560,V1232C1129,SI1232,end_vn1232);
V1233:VNPU3_3 port map (start_vn,clk,rst,Lc1233,C74V1233,C561V1233,C1130V1233,V1233C74,V1233C561,V1233C1130,SI1233,end_vn1233);
V1234:VNPU3_3 port map (start_vn,clk,rst,Lc1234,C75V1234,C562V1234,C1131V1234,V1234C75,V1234C562,V1234C1131,SI1234,end_vn1234);
V1235:VNPU3_3 port map (start_vn,clk,rst,Lc1235,C76V1235,C563V1235,C1132V1235,V1235C76,V1235C563,V1235C1132,SI1235,end_vn1235);
V1236:VNPU3_3 port map (start_vn,clk,rst,Lc1236,C77V1236,C564V1236,C1133V1236,V1236C77,V1236C564,V1236C1133,SI1236,end_vn1236);
V1237:VNPU3_3 port map (start_vn,clk,rst,Lc1237,C78V1237,C565V1237,C1134V1237,V1237C78,V1237C565,V1237C1134,SI1237,end_vn1237);
V1238:VNPU3_3 port map (start_vn,clk,rst,Lc1238,C79V1238,C566V1238,C1135V1238,V1238C79,V1238C566,V1238C1135,SI1238,end_vn1238);
V1239:VNPU3_3 port map (start_vn,clk,rst,Lc1239,C80V1239,C567V1239,C1136V1239,V1239C80,V1239C567,V1239C1136,SI1239,end_vn1239);
V1240:VNPU3_3 port map (start_vn,clk,rst,Lc1240,C81V1240,C568V1240,C1137V1240,V1240C81,V1240C568,V1240C1137,SI1240,end_vn1240);
V1241:VNPU3_3 port map (start_vn,clk,rst,Lc1241,C82V1241,C569V1241,C1138V1241,V1241C82,V1241C569,V1241C1138,SI1241,end_vn1241);
V1242:VNPU3_3 port map (start_vn,clk,rst,Lc1242,C83V1242,C570V1242,C1139V1242,V1242C83,V1242C570,V1242C1139,SI1242,end_vn1242);
V1243:VNPU3_3 port map (start_vn,clk,rst,Lc1243,C84V1243,C571V1243,C1140V1243,V1243C84,V1243C571,V1243C1140,SI1243,end_vn1243);
V1244:VNPU3_3 port map (start_vn,clk,rst,Lc1244,C85V1244,C572V1244,C1141V1244,V1244C85,V1244C572,V1244C1141,SI1244,end_vn1244);
V1245:VNPU3_3 port map (start_vn,clk,rst,Lc1245,C86V1245,C573V1245,C1142V1245,V1245C86,V1245C573,V1245C1142,SI1245,end_vn1245);
V1246:VNPU3_3 port map (start_vn,clk,rst,Lc1246,C87V1246,C574V1246,C1143V1246,V1246C87,V1246C574,V1246C1143,SI1246,end_vn1246);
V1247:VNPU3_3 port map (start_vn,clk,rst,Lc1247,C88V1247,C575V1247,C1144V1247,V1247C88,V1247C575,V1247C1144,SI1247,end_vn1247);
V1248:VNPU3_3 port map (start_vn,clk,rst,Lc1248,C89V1248,C576V1248,C1145V1248,V1248C89,V1248C576,V1248C1145,SI1248,end_vn1248);
V1249:VNPU2_2 port map (start_vn,clk,rst,Lc1249,C1V1249,C97V1249,V1249C1,V1249C97,SI1249,end_vn1249);
V1250:VNPU2_2 port map (start_vn,clk,rst,Lc1250,C2V1250,C98V1250,V1250C2,V1250C98,SI1250,end_vn1250);
V1251:VNPU2_2 port map (start_vn,clk,rst,Lc1251,C3V1251,C99V1251,V1251C3,V1251C99,SI1251,end_vn1251);
V1252:VNPU2_2 port map (start_vn,clk,rst,Lc1252,C4V1252,C100V1252,V1252C4,V1252C100,SI1252,end_vn1252);
V1253:VNPU2_2 port map (start_vn,clk,rst,Lc1253,C5V1253,C101V1253,V1253C5,V1253C101,SI1253,end_vn1253);
V1254:VNPU2_2 port map (start_vn,clk,rst,Lc1254,C6V1254,C102V1254,V1254C6,V1254C102,SI1254,end_vn1254);
V1255:VNPU2_2 port map (start_vn,clk,rst,Lc1255,C7V1255,C103V1255,V1255C7,V1255C103,SI1255,end_vn1255);
V1256:VNPU2_2 port map (start_vn,clk,rst,Lc1256,C8V1256,C104V1256,V1256C8,V1256C104,SI1256,end_vn1256);
V1257:VNPU2_2 port map (start_vn,clk,rst,Lc1257,C9V1257,C105V1257,V1257C9,V1257C105,SI1257,end_vn1257);
V1258:VNPU2_2 port map (start_vn,clk,rst,Lc1258,C10V1258,C106V1258,V1258C10,V1258C106,SI1258,end_vn1258);
V1259:VNPU2_2 port map (start_vn,clk,rst,Lc1259,C11V1259,C107V1259,V1259C11,V1259C107,SI1259,end_vn1259);
V1260:VNPU2_2 port map (start_vn,clk,rst,Lc1260,C12V1260,C108V1260,V1260C12,V1260C108,SI1260,end_vn1260);
V1261:VNPU2_2 port map (start_vn,clk,rst,Lc1261,C13V1261,C109V1261,V1261C13,V1261C109,SI1261,end_vn1261);
V1262:VNPU2_2 port map (start_vn,clk,rst,Lc1262,C14V1262,C110V1262,V1262C14,V1262C110,SI1262,end_vn1262);
V1263:VNPU2_2 port map (start_vn,clk,rst,Lc1263,C15V1263,C111V1263,V1263C15,V1263C111,SI1263,end_vn1263);
V1264:VNPU2_2 port map (start_vn,clk,rst,Lc1264,C16V1264,C112V1264,V1264C16,V1264C112,SI1264,end_vn1264);
V1265:VNPU2_2 port map (start_vn,clk,rst,Lc1265,C17V1265,C113V1265,V1265C17,V1265C113,SI1265,end_vn1265);
V1266:VNPU2_2 port map (start_vn,clk,rst,Lc1266,C18V1266,C114V1266,V1266C18,V1266C114,SI1266,end_vn1266);
V1267:VNPU2_2 port map (start_vn,clk,rst,Lc1267,C19V1267,C115V1267,V1267C19,V1267C115,SI1267,end_vn1267);
V1268:VNPU2_2 port map (start_vn,clk,rst,Lc1268,C20V1268,C116V1268,V1268C20,V1268C116,SI1268,end_vn1268);
V1269:VNPU2_2 port map (start_vn,clk,rst,Lc1269,C21V1269,C117V1269,V1269C21,V1269C117,SI1269,end_vn1269);
V1270:VNPU2_2 port map (start_vn,clk,rst,Lc1270,C22V1270,C118V1270,V1270C22,V1270C118,SI1270,end_vn1270);
V1271:VNPU2_2 port map (start_vn,clk,rst,Lc1271,C23V1271,C119V1271,V1271C23,V1271C119,SI1271,end_vn1271);
V1272:VNPU2_2 port map (start_vn,clk,rst,Lc1272,C24V1272,C120V1272,V1272C24,V1272C120,SI1272,end_vn1272);
V1273:VNPU2_2 port map (start_vn,clk,rst,Lc1273,C25V1273,C121V1273,V1273C25,V1273C121,SI1273,end_vn1273);
V1274:VNPU2_2 port map (start_vn,clk,rst,Lc1274,C26V1274,C122V1274,V1274C26,V1274C122,SI1274,end_vn1274);
V1275:VNPU2_2 port map (start_vn,clk,rst,Lc1275,C27V1275,C123V1275,V1275C27,V1275C123,SI1275,end_vn1275);
V1276:VNPU2_2 port map (start_vn,clk,rst,Lc1276,C28V1276,C124V1276,V1276C28,V1276C124,SI1276,end_vn1276);
V1277:VNPU2_2 port map (start_vn,clk,rst,Lc1277,C29V1277,C125V1277,V1277C29,V1277C125,SI1277,end_vn1277);
V1278:VNPU2_2 port map (start_vn,clk,rst,Lc1278,C30V1278,C126V1278,V1278C30,V1278C126,SI1278,end_vn1278);
V1279:VNPU2_2 port map (start_vn,clk,rst,Lc1279,C31V1279,C127V1279,V1279C31,V1279C127,SI1279,end_vn1279);
V1280:VNPU2_2 port map (start_vn,clk,rst,Lc1280,C32V1280,C128V1280,V1280C32,V1280C128,SI1280,end_vn1280);
V1281:VNPU2_2 port map (start_vn,clk,rst,Lc1281,C33V1281,C129V1281,V1281C33,V1281C129,SI1281,end_vn1281);
V1282:VNPU2_2 port map (start_vn,clk,rst,Lc1282,C34V1282,C130V1282,V1282C34,V1282C130,SI1282,end_vn1282);
V1283:VNPU2_2 port map (start_vn,clk,rst,Lc1283,C35V1283,C131V1283,V1283C35,V1283C131,SI1283,end_vn1283);
V1284:VNPU2_2 port map (start_vn,clk,rst,Lc1284,C36V1284,C132V1284,V1284C36,V1284C132,SI1284,end_vn1284);
V1285:VNPU2_2 port map (start_vn,clk,rst,Lc1285,C37V1285,C133V1285,V1285C37,V1285C133,SI1285,end_vn1285);
V1286:VNPU2_2 port map (start_vn,clk,rst,Lc1286,C38V1286,C134V1286,V1286C38,V1286C134,SI1286,end_vn1286);
V1287:VNPU2_2 port map (start_vn,clk,rst,Lc1287,C39V1287,C135V1287,V1287C39,V1287C135,SI1287,end_vn1287);
V1288:VNPU2_2 port map (start_vn,clk,rst,Lc1288,C40V1288,C136V1288,V1288C40,V1288C136,SI1288,end_vn1288);
V1289:VNPU2_2 port map (start_vn,clk,rst,Lc1289,C41V1289,C137V1289,V1289C41,V1289C137,SI1289,end_vn1289);
V1290:VNPU2_2 port map (start_vn,clk,rst,Lc1290,C42V1290,C138V1290,V1290C42,V1290C138,SI1290,end_vn1290);
V1291:VNPU2_2 port map (start_vn,clk,rst,Lc1291,C43V1291,C139V1291,V1291C43,V1291C139,SI1291,end_vn1291);
V1292:VNPU2_2 port map (start_vn,clk,rst,Lc1292,C44V1292,C140V1292,V1292C44,V1292C140,SI1292,end_vn1292);
V1293:VNPU2_2 port map (start_vn,clk,rst,Lc1293,C45V1293,C141V1293,V1293C45,V1293C141,SI1293,end_vn1293);
V1294:VNPU2_2 port map (start_vn,clk,rst,Lc1294,C46V1294,C142V1294,V1294C46,V1294C142,SI1294,end_vn1294);
V1295:VNPU2_2 port map (start_vn,clk,rst,Lc1295,C47V1295,C143V1295,V1295C47,V1295C143,SI1295,end_vn1295);
V1296:VNPU2_2 port map (start_vn,clk,rst,Lc1296,C48V1296,C144V1296,V1296C48,V1296C144,SI1296,end_vn1296);
V1297:VNPU2_2 port map (start_vn,clk,rst,Lc1297,C49V1297,C145V1297,V1297C49,V1297C145,SI1297,end_vn1297);
V1298:VNPU2_2 port map (start_vn,clk,rst,Lc1298,C50V1298,C146V1298,V1298C50,V1298C146,SI1298,end_vn1298);
V1299:VNPU2_2 port map (start_vn,clk,rst,Lc1299,C51V1299,C147V1299,V1299C51,V1299C147,SI1299,end_vn1299);
V1300:VNPU2_2 port map (start_vn,clk,rst,Lc1300,C52V1300,C148V1300,V1300C52,V1300C148,SI1300,end_vn1300);
V1301:VNPU2_2 port map (start_vn,clk,rst,Lc1301,C53V1301,C149V1301,V1301C53,V1301C149,SI1301,end_vn1301);
V1302:VNPU2_2 port map (start_vn,clk,rst,Lc1302,C54V1302,C150V1302,V1302C54,V1302C150,SI1302,end_vn1302);
V1303:VNPU2_2 port map (start_vn,clk,rst,Lc1303,C55V1303,C151V1303,V1303C55,V1303C151,SI1303,end_vn1303);
V1304:VNPU2_2 port map (start_vn,clk,rst,Lc1304,C56V1304,C152V1304,V1304C56,V1304C152,SI1304,end_vn1304);
V1305:VNPU2_2 port map (start_vn,clk,rst,Lc1305,C57V1305,C153V1305,V1305C57,V1305C153,SI1305,end_vn1305);
V1306:VNPU2_2 port map (start_vn,clk,rst,Lc1306,C58V1306,C154V1306,V1306C58,V1306C154,SI1306,end_vn1306);
V1307:VNPU2_2 port map (start_vn,clk,rst,Lc1307,C59V1307,C155V1307,V1307C59,V1307C155,SI1307,end_vn1307);
V1308:VNPU2_2 port map (start_vn,clk,rst,Lc1308,C60V1308,C156V1308,V1308C60,V1308C156,SI1308,end_vn1308);
V1309:VNPU2_2 port map (start_vn,clk,rst,Lc1309,C61V1309,C157V1309,V1309C61,V1309C157,SI1309,end_vn1309);
V1310:VNPU2_2 port map (start_vn,clk,rst,Lc1310,C62V1310,C158V1310,V1310C62,V1310C158,SI1310,end_vn1310);
V1311:VNPU2_2 port map (start_vn,clk,rst,Lc1311,C63V1311,C159V1311,V1311C63,V1311C159,SI1311,end_vn1311);
V1312:VNPU2_2 port map (start_vn,clk,rst,Lc1312,C64V1312,C160V1312,V1312C64,V1312C160,SI1312,end_vn1312);
V1313:VNPU2_2 port map (start_vn,clk,rst,Lc1313,C65V1313,C161V1313,V1313C65,V1313C161,SI1313,end_vn1313);
V1314:VNPU2_2 port map (start_vn,clk,rst,Lc1314,C66V1314,C162V1314,V1314C66,V1314C162,SI1314,end_vn1314);
V1315:VNPU2_2 port map (start_vn,clk,rst,Lc1315,C67V1315,C163V1315,V1315C67,V1315C163,SI1315,end_vn1315);
V1316:VNPU2_2 port map (start_vn,clk,rst,Lc1316,C68V1316,C164V1316,V1316C68,V1316C164,SI1316,end_vn1316);
V1317:VNPU2_2 port map (start_vn,clk,rst,Lc1317,C69V1317,C165V1317,V1317C69,V1317C165,SI1317,end_vn1317);
V1318:VNPU2_2 port map (start_vn,clk,rst,Lc1318,C70V1318,C166V1318,V1318C70,V1318C166,SI1318,end_vn1318);
V1319:VNPU2_2 port map (start_vn,clk,rst,Lc1319,C71V1319,C167V1319,V1319C71,V1319C167,SI1319,end_vn1319);
V1320:VNPU2_2 port map (start_vn,clk,rst,Lc1320,C72V1320,C168V1320,V1320C72,V1320C168,SI1320,end_vn1320);
V1321:VNPU2_2 port map (start_vn,clk,rst,Lc1321,C73V1321,C169V1321,V1321C73,V1321C169,SI1321,end_vn1321);
V1322:VNPU2_2 port map (start_vn,clk,rst,Lc1322,C74V1322,C170V1322,V1322C74,V1322C170,SI1322,end_vn1322);
V1323:VNPU2_2 port map (start_vn,clk,rst,Lc1323,C75V1323,C171V1323,V1323C75,V1323C171,SI1323,end_vn1323);
V1324:VNPU2_2 port map (start_vn,clk,rst,Lc1324,C76V1324,C172V1324,V1324C76,V1324C172,SI1324,end_vn1324);
V1325:VNPU2_2 port map (start_vn,clk,rst,Lc1325,C77V1325,C173V1325,V1325C77,V1325C173,SI1325,end_vn1325);
V1326:VNPU2_2 port map (start_vn,clk,rst,Lc1326,C78V1326,C174V1326,V1326C78,V1326C174,SI1326,end_vn1326);
V1327:VNPU2_2 port map (start_vn,clk,rst,Lc1327,C79V1327,C175V1327,V1327C79,V1327C175,SI1327,end_vn1327);
V1328:VNPU2_2 port map (start_vn,clk,rst,Lc1328,C80V1328,C176V1328,V1328C80,V1328C176,SI1328,end_vn1328);
V1329:VNPU2_2 port map (start_vn,clk,rst,Lc1329,C81V1329,C177V1329,V1329C81,V1329C177,SI1329,end_vn1329);
V1330:VNPU2_2 port map (start_vn,clk,rst,Lc1330,C82V1330,C178V1330,V1330C82,V1330C178,SI1330,end_vn1330);
V1331:VNPU2_2 port map (start_vn,clk,rst,Lc1331,C83V1331,C179V1331,V1331C83,V1331C179,SI1331,end_vn1331);
V1332:VNPU2_2 port map (start_vn,clk,rst,Lc1332,C84V1332,C180V1332,V1332C84,V1332C180,SI1332,end_vn1332);
V1333:VNPU2_2 port map (start_vn,clk,rst,Lc1333,C85V1333,C181V1333,V1333C85,V1333C181,SI1333,end_vn1333);
V1334:VNPU2_2 port map (start_vn,clk,rst,Lc1334,C86V1334,C182V1334,V1334C86,V1334C182,SI1334,end_vn1334);
V1335:VNPU2_2 port map (start_vn,clk,rst,Lc1335,C87V1335,C183V1335,V1335C87,V1335C183,SI1335,end_vn1335);
V1336:VNPU2_2 port map (start_vn,clk,rst,Lc1336,C88V1336,C184V1336,V1336C88,V1336C184,SI1336,end_vn1336);
V1337:VNPU2_2 port map (start_vn,clk,rst,Lc1337,C89V1337,C185V1337,V1337C89,V1337C185,SI1337,end_vn1337);
V1338:VNPU2_2 port map (start_vn,clk,rst,Lc1338,C90V1338,C186V1338,V1338C90,V1338C186,SI1338,end_vn1338);
V1339:VNPU2_2 port map (start_vn,clk,rst,Lc1339,C91V1339,C187V1339,V1339C91,V1339C187,SI1339,end_vn1339);
V1340:VNPU2_2 port map (start_vn,clk,rst,Lc1340,C92V1340,C188V1340,V1340C92,V1340C188,SI1340,end_vn1340);
V1341:VNPU2_2 port map (start_vn,clk,rst,Lc1341,C93V1341,C189V1341,V1341C93,V1341C189,SI1341,end_vn1341);
V1342:VNPU2_2 port map (start_vn,clk,rst,Lc1342,C94V1342,C190V1342,V1342C94,V1342C190,SI1342,end_vn1342);
V1343:VNPU2_2 port map (start_vn,clk,rst,Lc1343,C95V1343,C191V1343,V1343C95,V1343C191,SI1343,end_vn1343);
V1344:VNPU2_2 port map (start_vn,clk,rst,Lc1344,C96V1344,C192V1344,V1344C96,V1344C192,SI1344,end_vn1344);
V1345:VNPU2_2 port map (start_vn,clk,rst,Lc1345,C97V1345,C193V1345,V1345C97,V1345C193,SI1345,end_vn1345);
V1346:VNPU2_2 port map (start_vn,clk,rst,Lc1346,C98V1346,C194V1346,V1346C98,V1346C194,SI1346,end_vn1346);
V1347:VNPU2_2 port map (start_vn,clk,rst,Lc1347,C99V1347,C195V1347,V1347C99,V1347C195,SI1347,end_vn1347);
V1348:VNPU2_2 port map (start_vn,clk,rst,Lc1348,C100V1348,C196V1348,V1348C100,V1348C196,SI1348,end_vn1348);
V1349:VNPU2_2 port map (start_vn,clk,rst,Lc1349,C101V1349,C197V1349,V1349C101,V1349C197,SI1349,end_vn1349);
V1350:VNPU2_2 port map (start_vn,clk,rst,Lc1350,C102V1350,C198V1350,V1350C102,V1350C198,SI1350,end_vn1350);
V1351:VNPU2_2 port map (start_vn,clk,rst,Lc1351,C103V1351,C199V1351,V1351C103,V1351C199,SI1351,end_vn1351);
V1352:VNPU2_2 port map (start_vn,clk,rst,Lc1352,C104V1352,C200V1352,V1352C104,V1352C200,SI1352,end_vn1352);
V1353:VNPU2_2 port map (start_vn,clk,rst,Lc1353,C105V1353,C201V1353,V1353C105,V1353C201,SI1353,end_vn1353);
V1354:VNPU2_2 port map (start_vn,clk,rst,Lc1354,C106V1354,C202V1354,V1354C106,V1354C202,SI1354,end_vn1354);
V1355:VNPU2_2 port map (start_vn,clk,rst,Lc1355,C107V1355,C203V1355,V1355C107,V1355C203,SI1355,end_vn1355);
V1356:VNPU2_2 port map (start_vn,clk,rst,Lc1356,C108V1356,C204V1356,V1356C108,V1356C204,SI1356,end_vn1356);
V1357:VNPU2_2 port map (start_vn,clk,rst,Lc1357,C109V1357,C205V1357,V1357C109,V1357C205,SI1357,end_vn1357);
V1358:VNPU2_2 port map (start_vn,clk,rst,Lc1358,C110V1358,C206V1358,V1358C110,V1358C206,SI1358,end_vn1358);
V1359:VNPU2_2 port map (start_vn,clk,rst,Lc1359,C111V1359,C207V1359,V1359C111,V1359C207,SI1359,end_vn1359);
V1360:VNPU2_2 port map (start_vn,clk,rst,Lc1360,C112V1360,C208V1360,V1360C112,V1360C208,SI1360,end_vn1360);
V1361:VNPU2_2 port map (start_vn,clk,rst,Lc1361,C113V1361,C209V1361,V1361C113,V1361C209,SI1361,end_vn1361);
V1362:VNPU2_2 port map (start_vn,clk,rst,Lc1362,C114V1362,C210V1362,V1362C114,V1362C210,SI1362,end_vn1362);
V1363:VNPU2_2 port map (start_vn,clk,rst,Lc1363,C115V1363,C211V1363,V1363C115,V1363C211,SI1363,end_vn1363);
V1364:VNPU2_2 port map (start_vn,clk,rst,Lc1364,C116V1364,C212V1364,V1364C116,V1364C212,SI1364,end_vn1364);
V1365:VNPU2_2 port map (start_vn,clk,rst,Lc1365,C117V1365,C213V1365,V1365C117,V1365C213,SI1365,end_vn1365);
V1366:VNPU2_2 port map (start_vn,clk,rst,Lc1366,C118V1366,C214V1366,V1366C118,V1366C214,SI1366,end_vn1366);
V1367:VNPU2_2 port map (start_vn,clk,rst,Lc1367,C119V1367,C215V1367,V1367C119,V1367C215,SI1367,end_vn1367);
V1368:VNPU2_2 port map (start_vn,clk,rst,Lc1368,C120V1368,C216V1368,V1368C120,V1368C216,SI1368,end_vn1368);
V1369:VNPU2_2 port map (start_vn,clk,rst,Lc1369,C121V1369,C217V1369,V1369C121,V1369C217,SI1369,end_vn1369);
V1370:VNPU2_2 port map (start_vn,clk,rst,Lc1370,C122V1370,C218V1370,V1370C122,V1370C218,SI1370,end_vn1370);
V1371:VNPU2_2 port map (start_vn,clk,rst,Lc1371,C123V1371,C219V1371,V1371C123,V1371C219,SI1371,end_vn1371);
V1372:VNPU2_2 port map (start_vn,clk,rst,Lc1372,C124V1372,C220V1372,V1372C124,V1372C220,SI1372,end_vn1372);
V1373:VNPU2_2 port map (start_vn,clk,rst,Lc1373,C125V1373,C221V1373,V1373C125,V1373C221,SI1373,end_vn1373);
V1374:VNPU2_2 port map (start_vn,clk,rst,Lc1374,C126V1374,C222V1374,V1374C126,V1374C222,SI1374,end_vn1374);
V1375:VNPU2_2 port map (start_vn,clk,rst,Lc1375,C127V1375,C223V1375,V1375C127,V1375C223,SI1375,end_vn1375);
V1376:VNPU2_2 port map (start_vn,clk,rst,Lc1376,C128V1376,C224V1376,V1376C128,V1376C224,SI1376,end_vn1376);
V1377:VNPU2_2 port map (start_vn,clk,rst,Lc1377,C129V1377,C225V1377,V1377C129,V1377C225,SI1377,end_vn1377);
V1378:VNPU2_2 port map (start_vn,clk,rst,Lc1378,C130V1378,C226V1378,V1378C130,V1378C226,SI1378,end_vn1378);
V1379:VNPU2_2 port map (start_vn,clk,rst,Lc1379,C131V1379,C227V1379,V1379C131,V1379C227,SI1379,end_vn1379);
V1380:VNPU2_2 port map (start_vn,clk,rst,Lc1380,C132V1380,C228V1380,V1380C132,V1380C228,SI1380,end_vn1380);
V1381:VNPU2_2 port map (start_vn,clk,rst,Lc1381,C133V1381,C229V1381,V1381C133,V1381C229,SI1381,end_vn1381);
V1382:VNPU2_2 port map (start_vn,clk,rst,Lc1382,C134V1382,C230V1382,V1382C134,V1382C230,SI1382,end_vn1382);
V1383:VNPU2_2 port map (start_vn,clk,rst,Lc1383,C135V1383,C231V1383,V1383C135,V1383C231,SI1383,end_vn1383);
V1384:VNPU2_2 port map (start_vn,clk,rst,Lc1384,C136V1384,C232V1384,V1384C136,V1384C232,SI1384,end_vn1384);
V1385:VNPU2_2 port map (start_vn,clk,rst,Lc1385,C137V1385,C233V1385,V1385C137,V1385C233,SI1385,end_vn1385);
V1386:VNPU2_2 port map (start_vn,clk,rst,Lc1386,C138V1386,C234V1386,V1386C138,V1386C234,SI1386,end_vn1386);
V1387:VNPU2_2 port map (start_vn,clk,rst,Lc1387,C139V1387,C235V1387,V1387C139,V1387C235,SI1387,end_vn1387);
V1388:VNPU2_2 port map (start_vn,clk,rst,Lc1388,C140V1388,C236V1388,V1388C140,V1388C236,SI1388,end_vn1388);
V1389:VNPU2_2 port map (start_vn,clk,rst,Lc1389,C141V1389,C237V1389,V1389C141,V1389C237,SI1389,end_vn1389);
V1390:VNPU2_2 port map (start_vn,clk,rst,Lc1390,C142V1390,C238V1390,V1390C142,V1390C238,SI1390,end_vn1390);
V1391:VNPU2_2 port map (start_vn,clk,rst,Lc1391,C143V1391,C239V1391,V1391C143,V1391C239,SI1391,end_vn1391);
V1392:VNPU2_2 port map (start_vn,clk,rst,Lc1392,C144V1392,C240V1392,V1392C144,V1392C240,SI1392,end_vn1392);
V1393:VNPU2_2 port map (start_vn,clk,rst,Lc1393,C145V1393,C241V1393,V1393C145,V1393C241,SI1393,end_vn1393);
V1394:VNPU2_2 port map (start_vn,clk,rst,Lc1394,C146V1394,C242V1394,V1394C146,V1394C242,SI1394,end_vn1394);
V1395:VNPU2_2 port map (start_vn,clk,rst,Lc1395,C147V1395,C243V1395,V1395C147,V1395C243,SI1395,end_vn1395);
V1396:VNPU2_2 port map (start_vn,clk,rst,Lc1396,C148V1396,C244V1396,V1396C148,V1396C244,SI1396,end_vn1396);
V1397:VNPU2_2 port map (start_vn,clk,rst,Lc1397,C149V1397,C245V1397,V1397C149,V1397C245,SI1397,end_vn1397);
V1398:VNPU2_2 port map (start_vn,clk,rst,Lc1398,C150V1398,C246V1398,V1398C150,V1398C246,SI1398,end_vn1398);
V1399:VNPU2_2 port map (start_vn,clk,rst,Lc1399,C151V1399,C247V1399,V1399C151,V1399C247,SI1399,end_vn1399);
V1400:VNPU2_2 port map (start_vn,clk,rst,Lc1400,C152V1400,C248V1400,V1400C152,V1400C248,SI1400,end_vn1400);
V1401:VNPU2_2 port map (start_vn,clk,rst,Lc1401,C153V1401,C249V1401,V1401C153,V1401C249,SI1401,end_vn1401);
V1402:VNPU2_2 port map (start_vn,clk,rst,Lc1402,C154V1402,C250V1402,V1402C154,V1402C250,SI1402,end_vn1402);
V1403:VNPU2_2 port map (start_vn,clk,rst,Lc1403,C155V1403,C251V1403,V1403C155,V1403C251,SI1403,end_vn1403);
V1404:VNPU2_2 port map (start_vn,clk,rst,Lc1404,C156V1404,C252V1404,V1404C156,V1404C252,SI1404,end_vn1404);
V1405:VNPU2_2 port map (start_vn,clk,rst,Lc1405,C157V1405,C253V1405,V1405C157,V1405C253,SI1405,end_vn1405);
V1406:VNPU2_2 port map (start_vn,clk,rst,Lc1406,C158V1406,C254V1406,V1406C158,V1406C254,SI1406,end_vn1406);
V1407:VNPU2_2 port map (start_vn,clk,rst,Lc1407,C159V1407,C255V1407,V1407C159,V1407C255,SI1407,end_vn1407);
V1408:VNPU2_2 port map (start_vn,clk,rst,Lc1408,C160V1408,C256V1408,V1408C160,V1408C256,SI1408,end_vn1408);
V1409:VNPU2_2 port map (start_vn,clk,rst,Lc1409,C161V1409,C257V1409,V1409C161,V1409C257,SI1409,end_vn1409);
V1410:VNPU2_2 port map (start_vn,clk,rst,Lc1410,C162V1410,C258V1410,V1410C162,V1410C258,SI1410,end_vn1410);
V1411:VNPU2_2 port map (start_vn,clk,rst,Lc1411,C163V1411,C259V1411,V1411C163,V1411C259,SI1411,end_vn1411);
V1412:VNPU2_2 port map (start_vn,clk,rst,Lc1412,C164V1412,C260V1412,V1412C164,V1412C260,SI1412,end_vn1412);
V1413:VNPU2_2 port map (start_vn,clk,rst,Lc1413,C165V1413,C261V1413,V1413C165,V1413C261,SI1413,end_vn1413);
V1414:VNPU2_2 port map (start_vn,clk,rst,Lc1414,C166V1414,C262V1414,V1414C166,V1414C262,SI1414,end_vn1414);
V1415:VNPU2_2 port map (start_vn,clk,rst,Lc1415,C167V1415,C263V1415,V1415C167,V1415C263,SI1415,end_vn1415);
V1416:VNPU2_2 port map (start_vn,clk,rst,Lc1416,C168V1416,C264V1416,V1416C168,V1416C264,SI1416,end_vn1416);
V1417:VNPU2_2 port map (start_vn,clk,rst,Lc1417,C169V1417,C265V1417,V1417C169,V1417C265,SI1417,end_vn1417);
V1418:VNPU2_2 port map (start_vn,clk,rst,Lc1418,C170V1418,C266V1418,V1418C170,V1418C266,SI1418,end_vn1418);
V1419:VNPU2_2 port map (start_vn,clk,rst,Lc1419,C171V1419,C267V1419,V1419C171,V1419C267,SI1419,end_vn1419);
V1420:VNPU2_2 port map (start_vn,clk,rst,Lc1420,C172V1420,C268V1420,V1420C172,V1420C268,SI1420,end_vn1420);
V1421:VNPU2_2 port map (start_vn,clk,rst,Lc1421,C173V1421,C269V1421,V1421C173,V1421C269,SI1421,end_vn1421);
V1422:VNPU2_2 port map (start_vn,clk,rst,Lc1422,C174V1422,C270V1422,V1422C174,V1422C270,SI1422,end_vn1422);
V1423:VNPU2_2 port map (start_vn,clk,rst,Lc1423,C175V1423,C271V1423,V1423C175,V1423C271,SI1423,end_vn1423);
V1424:VNPU2_2 port map (start_vn,clk,rst,Lc1424,C176V1424,C272V1424,V1424C176,V1424C272,SI1424,end_vn1424);
V1425:VNPU2_2 port map (start_vn,clk,rst,Lc1425,C177V1425,C273V1425,V1425C177,V1425C273,SI1425,end_vn1425);
V1426:VNPU2_2 port map (start_vn,clk,rst,Lc1426,C178V1426,C274V1426,V1426C178,V1426C274,SI1426,end_vn1426);
V1427:VNPU2_2 port map (start_vn,clk,rst,Lc1427,C179V1427,C275V1427,V1427C179,V1427C275,SI1427,end_vn1427);
V1428:VNPU2_2 port map (start_vn,clk,rst,Lc1428,C180V1428,C276V1428,V1428C180,V1428C276,SI1428,end_vn1428);
V1429:VNPU2_2 port map (start_vn,clk,rst,Lc1429,C181V1429,C277V1429,V1429C181,V1429C277,SI1429,end_vn1429);
V1430:VNPU2_2 port map (start_vn,clk,rst,Lc1430,C182V1430,C278V1430,V1430C182,V1430C278,SI1430,end_vn1430);
V1431:VNPU2_2 port map (start_vn,clk,rst,Lc1431,C183V1431,C279V1431,V1431C183,V1431C279,SI1431,end_vn1431);
V1432:VNPU2_2 port map (start_vn,clk,rst,Lc1432,C184V1432,C280V1432,V1432C184,V1432C280,SI1432,end_vn1432);
V1433:VNPU2_2 port map (start_vn,clk,rst,Lc1433,C185V1433,C281V1433,V1433C185,V1433C281,SI1433,end_vn1433);
V1434:VNPU2_2 port map (start_vn,clk,rst,Lc1434,C186V1434,C282V1434,V1434C186,V1434C282,SI1434,end_vn1434);
V1435:VNPU2_2 port map (start_vn,clk,rst,Lc1435,C187V1435,C283V1435,V1435C187,V1435C283,SI1435,end_vn1435);
V1436:VNPU2_2 port map (start_vn,clk,rst,Lc1436,C188V1436,C284V1436,V1436C188,V1436C284,SI1436,end_vn1436);
V1437:VNPU2_2 port map (start_vn,clk,rst,Lc1437,C189V1437,C285V1437,V1437C189,V1437C285,SI1437,end_vn1437);
V1438:VNPU2_2 port map (start_vn,clk,rst,Lc1438,C190V1438,C286V1438,V1438C190,V1438C286,SI1438,end_vn1438);
V1439:VNPU2_2 port map (start_vn,clk,rst,Lc1439,C191V1439,C287V1439,V1439C191,V1439C287,SI1439,end_vn1439);
V1440:VNPU2_2 port map (start_vn,clk,rst,Lc1440,C192V1440,C288V1440,V1440C192,V1440C288,SI1440,end_vn1440);
V1441:VNPU2_2 port map (start_vn,clk,rst,Lc1441,C193V1441,C289V1441,V1441C193,V1441C289,SI1441,end_vn1441);
V1442:VNPU2_2 port map (start_vn,clk,rst,Lc1442,C194V1442,C290V1442,V1442C194,V1442C290,SI1442,end_vn1442);
V1443:VNPU2_2 port map (start_vn,clk,rst,Lc1443,C195V1443,C291V1443,V1443C195,V1443C291,SI1443,end_vn1443);
V1444:VNPU2_2 port map (start_vn,clk,rst,Lc1444,C196V1444,C292V1444,V1444C196,V1444C292,SI1444,end_vn1444);
V1445:VNPU2_2 port map (start_vn,clk,rst,Lc1445,C197V1445,C293V1445,V1445C197,V1445C293,SI1445,end_vn1445);
V1446:VNPU2_2 port map (start_vn,clk,rst,Lc1446,C198V1446,C294V1446,V1446C198,V1446C294,SI1446,end_vn1446);
V1447:VNPU2_2 port map (start_vn,clk,rst,Lc1447,C199V1447,C295V1447,V1447C199,V1447C295,SI1447,end_vn1447);
V1448:VNPU2_2 port map (start_vn,clk,rst,Lc1448,C200V1448,C296V1448,V1448C200,V1448C296,SI1448,end_vn1448);
V1449:VNPU2_2 port map (start_vn,clk,rst,Lc1449,C201V1449,C297V1449,V1449C201,V1449C297,SI1449,end_vn1449);
V1450:VNPU2_2 port map (start_vn,clk,rst,Lc1450,C202V1450,C298V1450,V1450C202,V1450C298,SI1450,end_vn1450);
V1451:VNPU2_2 port map (start_vn,clk,rst,Lc1451,C203V1451,C299V1451,V1451C203,V1451C299,SI1451,end_vn1451);
V1452:VNPU2_2 port map (start_vn,clk,rst,Lc1452,C204V1452,C300V1452,V1452C204,V1452C300,SI1452,end_vn1452);
V1453:VNPU2_2 port map (start_vn,clk,rst,Lc1453,C205V1453,C301V1453,V1453C205,V1453C301,SI1453,end_vn1453);
V1454:VNPU2_2 port map (start_vn,clk,rst,Lc1454,C206V1454,C302V1454,V1454C206,V1454C302,SI1454,end_vn1454);
V1455:VNPU2_2 port map (start_vn,clk,rst,Lc1455,C207V1455,C303V1455,V1455C207,V1455C303,SI1455,end_vn1455);
V1456:VNPU2_2 port map (start_vn,clk,rst,Lc1456,C208V1456,C304V1456,V1456C208,V1456C304,SI1456,end_vn1456);
V1457:VNPU2_2 port map (start_vn,clk,rst,Lc1457,C209V1457,C305V1457,V1457C209,V1457C305,SI1457,end_vn1457);
V1458:VNPU2_2 port map (start_vn,clk,rst,Lc1458,C210V1458,C306V1458,V1458C210,V1458C306,SI1458,end_vn1458);
V1459:VNPU2_2 port map (start_vn,clk,rst,Lc1459,C211V1459,C307V1459,V1459C211,V1459C307,SI1459,end_vn1459);
V1460:VNPU2_2 port map (start_vn,clk,rst,Lc1460,C212V1460,C308V1460,V1460C212,V1460C308,SI1460,end_vn1460);
V1461:VNPU2_2 port map (start_vn,clk,rst,Lc1461,C213V1461,C309V1461,V1461C213,V1461C309,SI1461,end_vn1461);
V1462:VNPU2_2 port map (start_vn,clk,rst,Lc1462,C214V1462,C310V1462,V1462C214,V1462C310,SI1462,end_vn1462);
V1463:VNPU2_2 port map (start_vn,clk,rst,Lc1463,C215V1463,C311V1463,V1463C215,V1463C311,SI1463,end_vn1463);
V1464:VNPU2_2 port map (start_vn,clk,rst,Lc1464,C216V1464,C312V1464,V1464C216,V1464C312,SI1464,end_vn1464);
V1465:VNPU2_2 port map (start_vn,clk,rst,Lc1465,C217V1465,C313V1465,V1465C217,V1465C313,SI1465,end_vn1465);
V1466:VNPU2_2 port map (start_vn,clk,rst,Lc1466,C218V1466,C314V1466,V1466C218,V1466C314,SI1466,end_vn1466);
V1467:VNPU2_2 port map (start_vn,clk,rst,Lc1467,C219V1467,C315V1467,V1467C219,V1467C315,SI1467,end_vn1467);
V1468:VNPU2_2 port map (start_vn,clk,rst,Lc1468,C220V1468,C316V1468,V1468C220,V1468C316,SI1468,end_vn1468);
V1469:VNPU2_2 port map (start_vn,clk,rst,Lc1469,C221V1469,C317V1469,V1469C221,V1469C317,SI1469,end_vn1469);
V1470:VNPU2_2 port map (start_vn,clk,rst,Lc1470,C222V1470,C318V1470,V1470C222,V1470C318,SI1470,end_vn1470);
V1471:VNPU2_2 port map (start_vn,clk,rst,Lc1471,C223V1471,C319V1471,V1471C223,V1471C319,SI1471,end_vn1471);
V1472:VNPU2_2 port map (start_vn,clk,rst,Lc1472,C224V1472,C320V1472,V1472C224,V1472C320,SI1472,end_vn1472);
V1473:VNPU2_2 port map (start_vn,clk,rst,Lc1473,C225V1473,C321V1473,V1473C225,V1473C321,SI1473,end_vn1473);
V1474:VNPU2_2 port map (start_vn,clk,rst,Lc1474,C226V1474,C322V1474,V1474C226,V1474C322,SI1474,end_vn1474);
V1475:VNPU2_2 port map (start_vn,clk,rst,Lc1475,C227V1475,C323V1475,V1475C227,V1475C323,SI1475,end_vn1475);
V1476:VNPU2_2 port map (start_vn,clk,rst,Lc1476,C228V1476,C324V1476,V1476C228,V1476C324,SI1476,end_vn1476);
V1477:VNPU2_2 port map (start_vn,clk,rst,Lc1477,C229V1477,C325V1477,V1477C229,V1477C325,SI1477,end_vn1477);
V1478:VNPU2_2 port map (start_vn,clk,rst,Lc1478,C230V1478,C326V1478,V1478C230,V1478C326,SI1478,end_vn1478);
V1479:VNPU2_2 port map (start_vn,clk,rst,Lc1479,C231V1479,C327V1479,V1479C231,V1479C327,SI1479,end_vn1479);
V1480:VNPU2_2 port map (start_vn,clk,rst,Lc1480,C232V1480,C328V1480,V1480C232,V1480C328,SI1480,end_vn1480);
V1481:VNPU2_2 port map (start_vn,clk,rst,Lc1481,C233V1481,C329V1481,V1481C233,V1481C329,SI1481,end_vn1481);
V1482:VNPU2_2 port map (start_vn,clk,rst,Lc1482,C234V1482,C330V1482,V1482C234,V1482C330,SI1482,end_vn1482);
V1483:VNPU2_2 port map (start_vn,clk,rst,Lc1483,C235V1483,C331V1483,V1483C235,V1483C331,SI1483,end_vn1483);
V1484:VNPU2_2 port map (start_vn,clk,rst,Lc1484,C236V1484,C332V1484,V1484C236,V1484C332,SI1484,end_vn1484);
V1485:VNPU2_2 port map (start_vn,clk,rst,Lc1485,C237V1485,C333V1485,V1485C237,V1485C333,SI1485,end_vn1485);
V1486:VNPU2_2 port map (start_vn,clk,rst,Lc1486,C238V1486,C334V1486,V1486C238,V1486C334,SI1486,end_vn1486);
V1487:VNPU2_2 port map (start_vn,clk,rst,Lc1487,C239V1487,C335V1487,V1487C239,V1487C335,SI1487,end_vn1487);
V1488:VNPU2_2 port map (start_vn,clk,rst,Lc1488,C240V1488,C336V1488,V1488C240,V1488C336,SI1488,end_vn1488);
V1489:VNPU2_2 port map (start_vn,clk,rst,Lc1489,C241V1489,C337V1489,V1489C241,V1489C337,SI1489,end_vn1489);
V1490:VNPU2_2 port map (start_vn,clk,rst,Lc1490,C242V1490,C338V1490,V1490C242,V1490C338,SI1490,end_vn1490);
V1491:VNPU2_2 port map (start_vn,clk,rst,Lc1491,C243V1491,C339V1491,V1491C243,V1491C339,SI1491,end_vn1491);
V1492:VNPU2_2 port map (start_vn,clk,rst,Lc1492,C244V1492,C340V1492,V1492C244,V1492C340,SI1492,end_vn1492);
V1493:VNPU2_2 port map (start_vn,clk,rst,Lc1493,C245V1493,C341V1493,V1493C245,V1493C341,SI1493,end_vn1493);
V1494:VNPU2_2 port map (start_vn,clk,rst,Lc1494,C246V1494,C342V1494,V1494C246,V1494C342,SI1494,end_vn1494);
V1495:VNPU2_2 port map (start_vn,clk,rst,Lc1495,C247V1495,C343V1495,V1495C247,V1495C343,SI1495,end_vn1495);
V1496:VNPU2_2 port map (start_vn,clk,rst,Lc1496,C248V1496,C344V1496,V1496C248,V1496C344,SI1496,end_vn1496);
V1497:VNPU2_2 port map (start_vn,clk,rst,Lc1497,C249V1497,C345V1497,V1497C249,V1497C345,SI1497,end_vn1497);
V1498:VNPU2_2 port map (start_vn,clk,rst,Lc1498,C250V1498,C346V1498,V1498C250,V1498C346,SI1498,end_vn1498);
V1499:VNPU2_2 port map (start_vn,clk,rst,Lc1499,C251V1499,C347V1499,V1499C251,V1499C347,SI1499,end_vn1499);
V1500:VNPU2_2 port map (start_vn,clk,rst,Lc1500,C252V1500,C348V1500,V1500C252,V1500C348,SI1500,end_vn1500);
V1501:VNPU2_2 port map (start_vn,clk,rst,Lc1501,C253V1501,C349V1501,V1501C253,V1501C349,SI1501,end_vn1501);
V1502:VNPU2_2 port map (start_vn,clk,rst,Lc1502,C254V1502,C350V1502,V1502C254,V1502C350,SI1502,end_vn1502);
V1503:VNPU2_2 port map (start_vn,clk,rst,Lc1503,C255V1503,C351V1503,V1503C255,V1503C351,SI1503,end_vn1503);
V1504:VNPU2_2 port map (start_vn,clk,rst,Lc1504,C256V1504,C352V1504,V1504C256,V1504C352,SI1504,end_vn1504);
V1505:VNPU2_2 port map (start_vn,clk,rst,Lc1505,C257V1505,C353V1505,V1505C257,V1505C353,SI1505,end_vn1505);
V1506:VNPU2_2 port map (start_vn,clk,rst,Lc1506,C258V1506,C354V1506,V1506C258,V1506C354,SI1506,end_vn1506);
V1507:VNPU2_2 port map (start_vn,clk,rst,Lc1507,C259V1507,C355V1507,V1507C259,V1507C355,SI1507,end_vn1507);
V1508:VNPU2_2 port map (start_vn,clk,rst,Lc1508,C260V1508,C356V1508,V1508C260,V1508C356,SI1508,end_vn1508);
V1509:VNPU2_2 port map (start_vn,clk,rst,Lc1509,C261V1509,C357V1509,V1509C261,V1509C357,SI1509,end_vn1509);
V1510:VNPU2_2 port map (start_vn,clk,rst,Lc1510,C262V1510,C358V1510,V1510C262,V1510C358,SI1510,end_vn1510);
V1511:VNPU2_2 port map (start_vn,clk,rst,Lc1511,C263V1511,C359V1511,V1511C263,V1511C359,SI1511,end_vn1511);
V1512:VNPU2_2 port map (start_vn,clk,rst,Lc1512,C264V1512,C360V1512,V1512C264,V1512C360,SI1512,end_vn1512);
V1513:VNPU2_2 port map (start_vn,clk,rst,Lc1513,C265V1513,C361V1513,V1513C265,V1513C361,SI1513,end_vn1513);
V1514:VNPU2_2 port map (start_vn,clk,rst,Lc1514,C266V1514,C362V1514,V1514C266,V1514C362,SI1514,end_vn1514);
V1515:VNPU2_2 port map (start_vn,clk,rst,Lc1515,C267V1515,C363V1515,V1515C267,V1515C363,SI1515,end_vn1515);
V1516:VNPU2_2 port map (start_vn,clk,rst,Lc1516,C268V1516,C364V1516,V1516C268,V1516C364,SI1516,end_vn1516);
V1517:VNPU2_2 port map (start_vn,clk,rst,Lc1517,C269V1517,C365V1517,V1517C269,V1517C365,SI1517,end_vn1517);
V1518:VNPU2_2 port map (start_vn,clk,rst,Lc1518,C270V1518,C366V1518,V1518C270,V1518C366,SI1518,end_vn1518);
V1519:VNPU2_2 port map (start_vn,clk,rst,Lc1519,C271V1519,C367V1519,V1519C271,V1519C367,SI1519,end_vn1519);
V1520:VNPU2_2 port map (start_vn,clk,rst,Lc1520,C272V1520,C368V1520,V1520C272,V1520C368,SI1520,end_vn1520);
V1521:VNPU2_2 port map (start_vn,clk,rst,Lc1521,C273V1521,C369V1521,V1521C273,V1521C369,SI1521,end_vn1521);
V1522:VNPU2_2 port map (start_vn,clk,rst,Lc1522,C274V1522,C370V1522,V1522C274,V1522C370,SI1522,end_vn1522);
V1523:VNPU2_2 port map (start_vn,clk,rst,Lc1523,C275V1523,C371V1523,V1523C275,V1523C371,SI1523,end_vn1523);
V1524:VNPU2_2 port map (start_vn,clk,rst,Lc1524,C276V1524,C372V1524,V1524C276,V1524C372,SI1524,end_vn1524);
V1525:VNPU2_2 port map (start_vn,clk,rst,Lc1525,C277V1525,C373V1525,V1525C277,V1525C373,SI1525,end_vn1525);
V1526:VNPU2_2 port map (start_vn,clk,rst,Lc1526,C278V1526,C374V1526,V1526C278,V1526C374,SI1526,end_vn1526);
V1527:VNPU2_2 port map (start_vn,clk,rst,Lc1527,C279V1527,C375V1527,V1527C279,V1527C375,SI1527,end_vn1527);
V1528:VNPU2_2 port map (start_vn,clk,rst,Lc1528,C280V1528,C376V1528,V1528C280,V1528C376,SI1528,end_vn1528);
V1529:VNPU2_2 port map (start_vn,clk,rst,Lc1529,C281V1529,C377V1529,V1529C281,V1529C377,SI1529,end_vn1529);
V1530:VNPU2_2 port map (start_vn,clk,rst,Lc1530,C282V1530,C378V1530,V1530C282,V1530C378,SI1530,end_vn1530);
V1531:VNPU2_2 port map (start_vn,clk,rst,Lc1531,C283V1531,C379V1531,V1531C283,V1531C379,SI1531,end_vn1531);
V1532:VNPU2_2 port map (start_vn,clk,rst,Lc1532,C284V1532,C380V1532,V1532C284,V1532C380,SI1532,end_vn1532);
V1533:VNPU2_2 port map (start_vn,clk,rst,Lc1533,C285V1533,C381V1533,V1533C285,V1533C381,SI1533,end_vn1533);
V1534:VNPU2_2 port map (start_vn,clk,rst,Lc1534,C286V1534,C382V1534,V1534C286,V1534C382,SI1534,end_vn1534);
V1535:VNPU2_2 port map (start_vn,clk,rst,Lc1535,C287V1535,C383V1535,V1535C287,V1535C383,SI1535,end_vn1535);
V1536:VNPU2_2 port map (start_vn,clk,rst,Lc1536,C288V1536,C384V1536,V1536C288,V1536C384,SI1536,end_vn1536);
V1537:VNPU2_2 port map (start_vn,clk,rst,Lc1537,C289V1537,C385V1537,V1537C289,V1537C385,SI1537,end_vn1537);
V1538:VNPU2_2 port map (start_vn,clk,rst,Lc1538,C290V1538,C386V1538,V1538C290,V1538C386,SI1538,end_vn1538);
V1539:VNPU2_2 port map (start_vn,clk,rst,Lc1539,C291V1539,C387V1539,V1539C291,V1539C387,SI1539,end_vn1539);
V1540:VNPU2_2 port map (start_vn,clk,rst,Lc1540,C292V1540,C388V1540,V1540C292,V1540C388,SI1540,end_vn1540);
V1541:VNPU2_2 port map (start_vn,clk,rst,Lc1541,C293V1541,C389V1541,V1541C293,V1541C389,SI1541,end_vn1541);
V1542:VNPU2_2 port map (start_vn,clk,rst,Lc1542,C294V1542,C390V1542,V1542C294,V1542C390,SI1542,end_vn1542);
V1543:VNPU2_2 port map (start_vn,clk,rst,Lc1543,C295V1543,C391V1543,V1543C295,V1543C391,SI1543,end_vn1543);
V1544:VNPU2_2 port map (start_vn,clk,rst,Lc1544,C296V1544,C392V1544,V1544C296,V1544C392,SI1544,end_vn1544);
V1545:VNPU2_2 port map (start_vn,clk,rst,Lc1545,C297V1545,C393V1545,V1545C297,V1545C393,SI1545,end_vn1545);
V1546:VNPU2_2 port map (start_vn,clk,rst,Lc1546,C298V1546,C394V1546,V1546C298,V1546C394,SI1546,end_vn1546);
V1547:VNPU2_2 port map (start_vn,clk,rst,Lc1547,C299V1547,C395V1547,V1547C299,V1547C395,SI1547,end_vn1547);
V1548:VNPU2_2 port map (start_vn,clk,rst,Lc1548,C300V1548,C396V1548,V1548C300,V1548C396,SI1548,end_vn1548);
V1549:VNPU2_2 port map (start_vn,clk,rst,Lc1549,C301V1549,C397V1549,V1549C301,V1549C397,SI1549,end_vn1549);
V1550:VNPU2_2 port map (start_vn,clk,rst,Lc1550,C302V1550,C398V1550,V1550C302,V1550C398,SI1550,end_vn1550);
V1551:VNPU2_2 port map (start_vn,clk,rst,Lc1551,C303V1551,C399V1551,V1551C303,V1551C399,SI1551,end_vn1551);
V1552:VNPU2_2 port map (start_vn,clk,rst,Lc1552,C304V1552,C400V1552,V1552C304,V1552C400,SI1552,end_vn1552);
V1553:VNPU2_2 port map (start_vn,clk,rst,Lc1553,C305V1553,C401V1553,V1553C305,V1553C401,SI1553,end_vn1553);
V1554:VNPU2_2 port map (start_vn,clk,rst,Lc1554,C306V1554,C402V1554,V1554C306,V1554C402,SI1554,end_vn1554);
V1555:VNPU2_2 port map (start_vn,clk,rst,Lc1555,C307V1555,C403V1555,V1555C307,V1555C403,SI1555,end_vn1555);
V1556:VNPU2_2 port map (start_vn,clk,rst,Lc1556,C308V1556,C404V1556,V1556C308,V1556C404,SI1556,end_vn1556);
V1557:VNPU2_2 port map (start_vn,clk,rst,Lc1557,C309V1557,C405V1557,V1557C309,V1557C405,SI1557,end_vn1557);
V1558:VNPU2_2 port map (start_vn,clk,rst,Lc1558,C310V1558,C406V1558,V1558C310,V1558C406,SI1558,end_vn1558);
V1559:VNPU2_2 port map (start_vn,clk,rst,Lc1559,C311V1559,C407V1559,V1559C311,V1559C407,SI1559,end_vn1559);
V1560:VNPU2_2 port map (start_vn,clk,rst,Lc1560,C312V1560,C408V1560,V1560C312,V1560C408,SI1560,end_vn1560);
V1561:VNPU2_2 port map (start_vn,clk,rst,Lc1561,C313V1561,C409V1561,V1561C313,V1561C409,SI1561,end_vn1561);
V1562:VNPU2_2 port map (start_vn,clk,rst,Lc1562,C314V1562,C410V1562,V1562C314,V1562C410,SI1562,end_vn1562);
V1563:VNPU2_2 port map (start_vn,clk,rst,Lc1563,C315V1563,C411V1563,V1563C315,V1563C411,SI1563,end_vn1563);
V1564:VNPU2_2 port map (start_vn,clk,rst,Lc1564,C316V1564,C412V1564,V1564C316,V1564C412,SI1564,end_vn1564);
V1565:VNPU2_2 port map (start_vn,clk,rst,Lc1565,C317V1565,C413V1565,V1565C317,V1565C413,SI1565,end_vn1565);
V1566:VNPU2_2 port map (start_vn,clk,rst,Lc1566,C318V1566,C414V1566,V1566C318,V1566C414,SI1566,end_vn1566);
V1567:VNPU2_2 port map (start_vn,clk,rst,Lc1567,C319V1567,C415V1567,V1567C319,V1567C415,SI1567,end_vn1567);
V1568:VNPU2_2 port map (start_vn,clk,rst,Lc1568,C320V1568,C416V1568,V1568C320,V1568C416,SI1568,end_vn1568);
V1569:VNPU2_2 port map (start_vn,clk,rst,Lc1569,C321V1569,C417V1569,V1569C321,V1569C417,SI1569,end_vn1569);
V1570:VNPU2_2 port map (start_vn,clk,rst,Lc1570,C322V1570,C418V1570,V1570C322,V1570C418,SI1570,end_vn1570);
V1571:VNPU2_2 port map (start_vn,clk,rst,Lc1571,C323V1571,C419V1571,V1571C323,V1571C419,SI1571,end_vn1571);
V1572:VNPU2_2 port map (start_vn,clk,rst,Lc1572,C324V1572,C420V1572,V1572C324,V1572C420,SI1572,end_vn1572);
V1573:VNPU2_2 port map (start_vn,clk,rst,Lc1573,C325V1573,C421V1573,V1573C325,V1573C421,SI1573,end_vn1573);
V1574:VNPU2_2 port map (start_vn,clk,rst,Lc1574,C326V1574,C422V1574,V1574C326,V1574C422,SI1574,end_vn1574);
V1575:VNPU2_2 port map (start_vn,clk,rst,Lc1575,C327V1575,C423V1575,V1575C327,V1575C423,SI1575,end_vn1575);
V1576:VNPU2_2 port map (start_vn,clk,rst,Lc1576,C328V1576,C424V1576,V1576C328,V1576C424,SI1576,end_vn1576);
V1577:VNPU2_2 port map (start_vn,clk,rst,Lc1577,C329V1577,C425V1577,V1577C329,V1577C425,SI1577,end_vn1577);
V1578:VNPU2_2 port map (start_vn,clk,rst,Lc1578,C330V1578,C426V1578,V1578C330,V1578C426,SI1578,end_vn1578);
V1579:VNPU2_2 port map (start_vn,clk,rst,Lc1579,C331V1579,C427V1579,V1579C331,V1579C427,SI1579,end_vn1579);
V1580:VNPU2_2 port map (start_vn,clk,rst,Lc1580,C332V1580,C428V1580,V1580C332,V1580C428,SI1580,end_vn1580);
V1581:VNPU2_2 port map (start_vn,clk,rst,Lc1581,C333V1581,C429V1581,V1581C333,V1581C429,SI1581,end_vn1581);
V1582:VNPU2_2 port map (start_vn,clk,rst,Lc1582,C334V1582,C430V1582,V1582C334,V1582C430,SI1582,end_vn1582);
V1583:VNPU2_2 port map (start_vn,clk,rst,Lc1583,C335V1583,C431V1583,V1583C335,V1583C431,SI1583,end_vn1583);
V1584:VNPU2_2 port map (start_vn,clk,rst,Lc1584,C336V1584,C432V1584,V1584C336,V1584C432,SI1584,end_vn1584);
V1585:VNPU2_2 port map (start_vn,clk,rst,Lc1585,C337V1585,C433V1585,V1585C337,V1585C433,SI1585,end_vn1585);
V1586:VNPU2_2 port map (start_vn,clk,rst,Lc1586,C338V1586,C434V1586,V1586C338,V1586C434,SI1586,end_vn1586);
V1587:VNPU2_2 port map (start_vn,clk,rst,Lc1587,C339V1587,C435V1587,V1587C339,V1587C435,SI1587,end_vn1587);
V1588:VNPU2_2 port map (start_vn,clk,rst,Lc1588,C340V1588,C436V1588,V1588C340,V1588C436,SI1588,end_vn1588);
V1589:VNPU2_2 port map (start_vn,clk,rst,Lc1589,C341V1589,C437V1589,V1589C341,V1589C437,SI1589,end_vn1589);
V1590:VNPU2_2 port map (start_vn,clk,rst,Lc1590,C342V1590,C438V1590,V1590C342,V1590C438,SI1590,end_vn1590);
V1591:VNPU2_2 port map (start_vn,clk,rst,Lc1591,C343V1591,C439V1591,V1591C343,V1591C439,SI1591,end_vn1591);
V1592:VNPU2_2 port map (start_vn,clk,rst,Lc1592,C344V1592,C440V1592,V1592C344,V1592C440,SI1592,end_vn1592);
V1593:VNPU2_2 port map (start_vn,clk,rst,Lc1593,C345V1593,C441V1593,V1593C345,V1593C441,SI1593,end_vn1593);
V1594:VNPU2_2 port map (start_vn,clk,rst,Lc1594,C346V1594,C442V1594,V1594C346,V1594C442,SI1594,end_vn1594);
V1595:VNPU2_2 port map (start_vn,clk,rst,Lc1595,C347V1595,C443V1595,V1595C347,V1595C443,SI1595,end_vn1595);
V1596:VNPU2_2 port map (start_vn,clk,rst,Lc1596,C348V1596,C444V1596,V1596C348,V1596C444,SI1596,end_vn1596);
V1597:VNPU2_2 port map (start_vn,clk,rst,Lc1597,C349V1597,C445V1597,V1597C349,V1597C445,SI1597,end_vn1597);
V1598:VNPU2_2 port map (start_vn,clk,rst,Lc1598,C350V1598,C446V1598,V1598C350,V1598C446,SI1598,end_vn1598);
V1599:VNPU2_2 port map (start_vn,clk,rst,Lc1599,C351V1599,C447V1599,V1599C351,V1599C447,SI1599,end_vn1599);
V1600:VNPU2_2 port map (start_vn,clk,rst,Lc1600,C352V1600,C448V1600,V1600C352,V1600C448,SI1600,end_vn1600);
V1601:VNPU2_2 port map (start_vn,clk,rst,Lc1601,C353V1601,C449V1601,V1601C353,V1601C449,SI1601,end_vn1601);
V1602:VNPU2_2 port map (start_vn,clk,rst,Lc1602,C354V1602,C450V1602,V1602C354,V1602C450,SI1602,end_vn1602);
V1603:VNPU2_2 port map (start_vn,clk,rst,Lc1603,C355V1603,C451V1603,V1603C355,V1603C451,SI1603,end_vn1603);
V1604:VNPU2_2 port map (start_vn,clk,rst,Lc1604,C356V1604,C452V1604,V1604C356,V1604C452,SI1604,end_vn1604);
V1605:VNPU2_2 port map (start_vn,clk,rst,Lc1605,C357V1605,C453V1605,V1605C357,V1605C453,SI1605,end_vn1605);
V1606:VNPU2_2 port map (start_vn,clk,rst,Lc1606,C358V1606,C454V1606,V1606C358,V1606C454,SI1606,end_vn1606);
V1607:VNPU2_2 port map (start_vn,clk,rst,Lc1607,C359V1607,C455V1607,V1607C359,V1607C455,SI1607,end_vn1607);
V1608:VNPU2_2 port map (start_vn,clk,rst,Lc1608,C360V1608,C456V1608,V1608C360,V1608C456,SI1608,end_vn1608);
V1609:VNPU2_2 port map (start_vn,clk,rst,Lc1609,C361V1609,C457V1609,V1609C361,V1609C457,SI1609,end_vn1609);
V1610:VNPU2_2 port map (start_vn,clk,rst,Lc1610,C362V1610,C458V1610,V1610C362,V1610C458,SI1610,end_vn1610);
V1611:VNPU2_2 port map (start_vn,clk,rst,Lc1611,C363V1611,C459V1611,V1611C363,V1611C459,SI1611,end_vn1611);
V1612:VNPU2_2 port map (start_vn,clk,rst,Lc1612,C364V1612,C460V1612,V1612C364,V1612C460,SI1612,end_vn1612);
V1613:VNPU2_2 port map (start_vn,clk,rst,Lc1613,C365V1613,C461V1613,V1613C365,V1613C461,SI1613,end_vn1613);
V1614:VNPU2_2 port map (start_vn,clk,rst,Lc1614,C366V1614,C462V1614,V1614C366,V1614C462,SI1614,end_vn1614);
V1615:VNPU2_2 port map (start_vn,clk,rst,Lc1615,C367V1615,C463V1615,V1615C367,V1615C463,SI1615,end_vn1615);
V1616:VNPU2_2 port map (start_vn,clk,rst,Lc1616,C368V1616,C464V1616,V1616C368,V1616C464,SI1616,end_vn1616);
V1617:VNPU2_2 port map (start_vn,clk,rst,Lc1617,C369V1617,C465V1617,V1617C369,V1617C465,SI1617,end_vn1617);
V1618:VNPU2_2 port map (start_vn,clk,rst,Lc1618,C370V1618,C466V1618,V1618C370,V1618C466,SI1618,end_vn1618);
V1619:VNPU2_2 port map (start_vn,clk,rst,Lc1619,C371V1619,C467V1619,V1619C371,V1619C467,SI1619,end_vn1619);
V1620:VNPU2_2 port map (start_vn,clk,rst,Lc1620,C372V1620,C468V1620,V1620C372,V1620C468,SI1620,end_vn1620);
V1621:VNPU2_2 port map (start_vn,clk,rst,Lc1621,C373V1621,C469V1621,V1621C373,V1621C469,SI1621,end_vn1621);
V1622:VNPU2_2 port map (start_vn,clk,rst,Lc1622,C374V1622,C470V1622,V1622C374,V1622C470,SI1622,end_vn1622);
V1623:VNPU2_2 port map (start_vn,clk,rst,Lc1623,C375V1623,C471V1623,V1623C375,V1623C471,SI1623,end_vn1623);
V1624:VNPU2_2 port map (start_vn,clk,rst,Lc1624,C376V1624,C472V1624,V1624C376,V1624C472,SI1624,end_vn1624);
V1625:VNPU2_2 port map (start_vn,clk,rst,Lc1625,C377V1625,C473V1625,V1625C377,V1625C473,SI1625,end_vn1625);
V1626:VNPU2_2 port map (start_vn,clk,rst,Lc1626,C378V1626,C474V1626,V1626C378,V1626C474,SI1626,end_vn1626);
V1627:VNPU2_2 port map (start_vn,clk,rst,Lc1627,C379V1627,C475V1627,V1627C379,V1627C475,SI1627,end_vn1627);
V1628:VNPU2_2 port map (start_vn,clk,rst,Lc1628,C380V1628,C476V1628,V1628C380,V1628C476,SI1628,end_vn1628);
V1629:VNPU2_2 port map (start_vn,clk,rst,Lc1629,C381V1629,C477V1629,V1629C381,V1629C477,SI1629,end_vn1629);
V1630:VNPU2_2 port map (start_vn,clk,rst,Lc1630,C382V1630,C478V1630,V1630C382,V1630C478,SI1630,end_vn1630);
V1631:VNPU2_2 port map (start_vn,clk,rst,Lc1631,C383V1631,C479V1631,V1631C383,V1631C479,SI1631,end_vn1631);
V1632:VNPU2_2 port map (start_vn,clk,rst,Lc1632,C384V1632,C480V1632,V1632C384,V1632C480,SI1632,end_vn1632);
V1633:VNPU2_2 port map (start_vn,clk,rst,Lc1633,C385V1633,C481V1633,V1633C385,V1633C481,SI1633,end_vn1633);
V1634:VNPU2_2 port map (start_vn,clk,rst,Lc1634,C386V1634,C482V1634,V1634C386,V1634C482,SI1634,end_vn1634);
V1635:VNPU2_2 port map (start_vn,clk,rst,Lc1635,C387V1635,C483V1635,V1635C387,V1635C483,SI1635,end_vn1635);
V1636:VNPU2_2 port map (start_vn,clk,rst,Lc1636,C388V1636,C484V1636,V1636C388,V1636C484,SI1636,end_vn1636);
V1637:VNPU2_2 port map (start_vn,clk,rst,Lc1637,C389V1637,C485V1637,V1637C389,V1637C485,SI1637,end_vn1637);
V1638:VNPU2_2 port map (start_vn,clk,rst,Lc1638,C390V1638,C486V1638,V1638C390,V1638C486,SI1638,end_vn1638);
V1639:VNPU2_2 port map (start_vn,clk,rst,Lc1639,C391V1639,C487V1639,V1639C391,V1639C487,SI1639,end_vn1639);
V1640:VNPU2_2 port map (start_vn,clk,rst,Lc1640,C392V1640,C488V1640,V1640C392,V1640C488,SI1640,end_vn1640);
V1641:VNPU2_2 port map (start_vn,clk,rst,Lc1641,C393V1641,C489V1641,V1641C393,V1641C489,SI1641,end_vn1641);
V1642:VNPU2_2 port map (start_vn,clk,rst,Lc1642,C394V1642,C490V1642,V1642C394,V1642C490,SI1642,end_vn1642);
V1643:VNPU2_2 port map (start_vn,clk,rst,Lc1643,C395V1643,C491V1643,V1643C395,V1643C491,SI1643,end_vn1643);
V1644:VNPU2_2 port map (start_vn,clk,rst,Lc1644,C396V1644,C492V1644,V1644C396,V1644C492,SI1644,end_vn1644);
V1645:VNPU2_2 port map (start_vn,clk,rst,Lc1645,C397V1645,C493V1645,V1645C397,V1645C493,SI1645,end_vn1645);
V1646:VNPU2_2 port map (start_vn,clk,rst,Lc1646,C398V1646,C494V1646,V1646C398,V1646C494,SI1646,end_vn1646);
V1647:VNPU2_2 port map (start_vn,clk,rst,Lc1647,C399V1647,C495V1647,V1647C399,V1647C495,SI1647,end_vn1647);
V1648:VNPU2_2 port map (start_vn,clk,rst,Lc1648,C400V1648,C496V1648,V1648C400,V1648C496,SI1648,end_vn1648);
V1649:VNPU2_2 port map (start_vn,clk,rst,Lc1649,C401V1649,C497V1649,V1649C401,V1649C497,SI1649,end_vn1649);
V1650:VNPU2_2 port map (start_vn,clk,rst,Lc1650,C402V1650,C498V1650,V1650C402,V1650C498,SI1650,end_vn1650);
V1651:VNPU2_2 port map (start_vn,clk,rst,Lc1651,C403V1651,C499V1651,V1651C403,V1651C499,SI1651,end_vn1651);
V1652:VNPU2_2 port map (start_vn,clk,rst,Lc1652,C404V1652,C500V1652,V1652C404,V1652C500,SI1652,end_vn1652);
V1653:VNPU2_2 port map (start_vn,clk,rst,Lc1653,C405V1653,C501V1653,V1653C405,V1653C501,SI1653,end_vn1653);
V1654:VNPU2_2 port map (start_vn,clk,rst,Lc1654,C406V1654,C502V1654,V1654C406,V1654C502,SI1654,end_vn1654);
V1655:VNPU2_2 port map (start_vn,clk,rst,Lc1655,C407V1655,C503V1655,V1655C407,V1655C503,SI1655,end_vn1655);
V1656:VNPU2_2 port map (start_vn,clk,rst,Lc1656,C408V1656,C504V1656,V1656C408,V1656C504,SI1656,end_vn1656);
V1657:VNPU2_2 port map (start_vn,clk,rst,Lc1657,C409V1657,C505V1657,V1657C409,V1657C505,SI1657,end_vn1657);
V1658:VNPU2_2 port map (start_vn,clk,rst,Lc1658,C410V1658,C506V1658,V1658C410,V1658C506,SI1658,end_vn1658);
V1659:VNPU2_2 port map (start_vn,clk,rst,Lc1659,C411V1659,C507V1659,V1659C411,V1659C507,SI1659,end_vn1659);
V1660:VNPU2_2 port map (start_vn,clk,rst,Lc1660,C412V1660,C508V1660,V1660C412,V1660C508,SI1660,end_vn1660);
V1661:VNPU2_2 port map (start_vn,clk,rst,Lc1661,C413V1661,C509V1661,V1661C413,V1661C509,SI1661,end_vn1661);
V1662:VNPU2_2 port map (start_vn,clk,rst,Lc1662,C414V1662,C510V1662,V1662C414,V1662C510,SI1662,end_vn1662);
V1663:VNPU2_2 port map (start_vn,clk,rst,Lc1663,C415V1663,C511V1663,V1663C415,V1663C511,SI1663,end_vn1663);
V1664:VNPU2_2 port map (start_vn,clk,rst,Lc1664,C416V1664,C512V1664,V1664C416,V1664C512,SI1664,end_vn1664);
V1665:VNPU2_2 port map (start_vn,clk,rst,Lc1665,C417V1665,C513V1665,V1665C417,V1665C513,SI1665,end_vn1665);
V1666:VNPU2_2 port map (start_vn,clk,rst,Lc1666,C418V1666,C514V1666,V1666C418,V1666C514,SI1666,end_vn1666);
V1667:VNPU2_2 port map (start_vn,clk,rst,Lc1667,C419V1667,C515V1667,V1667C419,V1667C515,SI1667,end_vn1667);
V1668:VNPU2_2 port map (start_vn,clk,rst,Lc1668,C420V1668,C516V1668,V1668C420,V1668C516,SI1668,end_vn1668);
V1669:VNPU2_2 port map (start_vn,clk,rst,Lc1669,C421V1669,C517V1669,V1669C421,V1669C517,SI1669,end_vn1669);
V1670:VNPU2_2 port map (start_vn,clk,rst,Lc1670,C422V1670,C518V1670,V1670C422,V1670C518,SI1670,end_vn1670);
V1671:VNPU2_2 port map (start_vn,clk,rst,Lc1671,C423V1671,C519V1671,V1671C423,V1671C519,SI1671,end_vn1671);
V1672:VNPU2_2 port map (start_vn,clk,rst,Lc1672,C424V1672,C520V1672,V1672C424,V1672C520,SI1672,end_vn1672);
V1673:VNPU2_2 port map (start_vn,clk,rst,Lc1673,C425V1673,C521V1673,V1673C425,V1673C521,SI1673,end_vn1673);
V1674:VNPU2_2 port map (start_vn,clk,rst,Lc1674,C426V1674,C522V1674,V1674C426,V1674C522,SI1674,end_vn1674);
V1675:VNPU2_2 port map (start_vn,clk,rst,Lc1675,C427V1675,C523V1675,V1675C427,V1675C523,SI1675,end_vn1675);
V1676:VNPU2_2 port map (start_vn,clk,rst,Lc1676,C428V1676,C524V1676,V1676C428,V1676C524,SI1676,end_vn1676);
V1677:VNPU2_2 port map (start_vn,clk,rst,Lc1677,C429V1677,C525V1677,V1677C429,V1677C525,SI1677,end_vn1677);
V1678:VNPU2_2 port map (start_vn,clk,rst,Lc1678,C430V1678,C526V1678,V1678C430,V1678C526,SI1678,end_vn1678);
V1679:VNPU2_2 port map (start_vn,clk,rst,Lc1679,C431V1679,C527V1679,V1679C431,V1679C527,SI1679,end_vn1679);
V1680:VNPU2_2 port map (start_vn,clk,rst,Lc1680,C432V1680,C528V1680,V1680C432,V1680C528,SI1680,end_vn1680);
V1681:VNPU2_2 port map (start_vn,clk,rst,Lc1681,C433V1681,C529V1681,V1681C433,V1681C529,SI1681,end_vn1681);
V1682:VNPU2_2 port map (start_vn,clk,rst,Lc1682,C434V1682,C530V1682,V1682C434,V1682C530,SI1682,end_vn1682);
V1683:VNPU2_2 port map (start_vn,clk,rst,Lc1683,C435V1683,C531V1683,V1683C435,V1683C531,SI1683,end_vn1683);
V1684:VNPU2_2 port map (start_vn,clk,rst,Lc1684,C436V1684,C532V1684,V1684C436,V1684C532,SI1684,end_vn1684);
V1685:VNPU2_2 port map (start_vn,clk,rst,Lc1685,C437V1685,C533V1685,V1685C437,V1685C533,SI1685,end_vn1685);
V1686:VNPU2_2 port map (start_vn,clk,rst,Lc1686,C438V1686,C534V1686,V1686C438,V1686C534,SI1686,end_vn1686);
V1687:VNPU2_2 port map (start_vn,clk,rst,Lc1687,C439V1687,C535V1687,V1687C439,V1687C535,SI1687,end_vn1687);
V1688:VNPU2_2 port map (start_vn,clk,rst,Lc1688,C440V1688,C536V1688,V1688C440,V1688C536,SI1688,end_vn1688);
V1689:VNPU2_2 port map (start_vn,clk,rst,Lc1689,C441V1689,C537V1689,V1689C441,V1689C537,SI1689,end_vn1689);
V1690:VNPU2_2 port map (start_vn,clk,rst,Lc1690,C442V1690,C538V1690,V1690C442,V1690C538,SI1690,end_vn1690);
V1691:VNPU2_2 port map (start_vn,clk,rst,Lc1691,C443V1691,C539V1691,V1691C443,V1691C539,SI1691,end_vn1691);
V1692:VNPU2_2 port map (start_vn,clk,rst,Lc1692,C444V1692,C540V1692,V1692C444,V1692C540,SI1692,end_vn1692);
V1693:VNPU2_2 port map (start_vn,clk,rst,Lc1693,C445V1693,C541V1693,V1693C445,V1693C541,SI1693,end_vn1693);
V1694:VNPU2_2 port map (start_vn,clk,rst,Lc1694,C446V1694,C542V1694,V1694C446,V1694C542,SI1694,end_vn1694);
V1695:VNPU2_2 port map (start_vn,clk,rst,Lc1695,C447V1695,C543V1695,V1695C447,V1695C543,SI1695,end_vn1695);
V1696:VNPU2_2 port map (start_vn,clk,rst,Lc1696,C448V1696,C544V1696,V1696C448,V1696C544,SI1696,end_vn1696);
V1697:VNPU2_2 port map (start_vn,clk,rst,Lc1697,C449V1697,C545V1697,V1697C449,V1697C545,SI1697,end_vn1697);
V1698:VNPU2_2 port map (start_vn,clk,rst,Lc1698,C450V1698,C546V1698,V1698C450,V1698C546,SI1698,end_vn1698);
V1699:VNPU2_2 port map (start_vn,clk,rst,Lc1699,C451V1699,C547V1699,V1699C451,V1699C547,SI1699,end_vn1699);
V1700:VNPU2_2 port map (start_vn,clk,rst,Lc1700,C452V1700,C548V1700,V1700C452,V1700C548,SI1700,end_vn1700);
V1701:VNPU2_2 port map (start_vn,clk,rst,Lc1701,C453V1701,C549V1701,V1701C453,V1701C549,SI1701,end_vn1701);
V1702:VNPU2_2 port map (start_vn,clk,rst,Lc1702,C454V1702,C550V1702,V1702C454,V1702C550,SI1702,end_vn1702);
V1703:VNPU2_2 port map (start_vn,clk,rst,Lc1703,C455V1703,C551V1703,V1703C455,V1703C551,SI1703,end_vn1703);
V1704:VNPU2_2 port map (start_vn,clk,rst,Lc1704,C456V1704,C552V1704,V1704C456,V1704C552,SI1704,end_vn1704);
V1705:VNPU2_2 port map (start_vn,clk,rst,Lc1705,C457V1705,C553V1705,V1705C457,V1705C553,SI1705,end_vn1705);
V1706:VNPU2_2 port map (start_vn,clk,rst,Lc1706,C458V1706,C554V1706,V1706C458,V1706C554,SI1706,end_vn1706);
V1707:VNPU2_2 port map (start_vn,clk,rst,Lc1707,C459V1707,C555V1707,V1707C459,V1707C555,SI1707,end_vn1707);
V1708:VNPU2_2 port map (start_vn,clk,rst,Lc1708,C460V1708,C556V1708,V1708C460,V1708C556,SI1708,end_vn1708);
V1709:VNPU2_2 port map (start_vn,clk,rst,Lc1709,C461V1709,C557V1709,V1709C461,V1709C557,SI1709,end_vn1709);
V1710:VNPU2_2 port map (start_vn,clk,rst,Lc1710,C462V1710,C558V1710,V1710C462,V1710C558,SI1710,end_vn1710);
V1711:VNPU2_2 port map (start_vn,clk,rst,Lc1711,C463V1711,C559V1711,V1711C463,V1711C559,SI1711,end_vn1711);
V1712:VNPU2_2 port map (start_vn,clk,rst,Lc1712,C464V1712,C560V1712,V1712C464,V1712C560,SI1712,end_vn1712);
V1713:VNPU2_2 port map (start_vn,clk,rst,Lc1713,C465V1713,C561V1713,V1713C465,V1713C561,SI1713,end_vn1713);
V1714:VNPU2_2 port map (start_vn,clk,rst,Lc1714,C466V1714,C562V1714,V1714C466,V1714C562,SI1714,end_vn1714);
V1715:VNPU2_2 port map (start_vn,clk,rst,Lc1715,C467V1715,C563V1715,V1715C467,V1715C563,SI1715,end_vn1715);
V1716:VNPU2_2 port map (start_vn,clk,rst,Lc1716,C468V1716,C564V1716,V1716C468,V1716C564,SI1716,end_vn1716);
V1717:VNPU2_2 port map (start_vn,clk,rst,Lc1717,C469V1717,C565V1717,V1717C469,V1717C565,SI1717,end_vn1717);
V1718:VNPU2_2 port map (start_vn,clk,rst,Lc1718,C470V1718,C566V1718,V1718C470,V1718C566,SI1718,end_vn1718);
V1719:VNPU2_2 port map (start_vn,clk,rst,Lc1719,C471V1719,C567V1719,V1719C471,V1719C567,SI1719,end_vn1719);
V1720:VNPU2_2 port map (start_vn,clk,rst,Lc1720,C472V1720,C568V1720,V1720C472,V1720C568,SI1720,end_vn1720);
V1721:VNPU2_2 port map (start_vn,clk,rst,Lc1721,C473V1721,C569V1721,V1721C473,V1721C569,SI1721,end_vn1721);
V1722:VNPU2_2 port map (start_vn,clk,rst,Lc1722,C474V1722,C570V1722,V1722C474,V1722C570,SI1722,end_vn1722);
V1723:VNPU2_2 port map (start_vn,clk,rst,Lc1723,C475V1723,C571V1723,V1723C475,V1723C571,SI1723,end_vn1723);
V1724:VNPU2_2 port map (start_vn,clk,rst,Lc1724,C476V1724,C572V1724,V1724C476,V1724C572,SI1724,end_vn1724);
V1725:VNPU2_2 port map (start_vn,clk,rst,Lc1725,C477V1725,C573V1725,V1725C477,V1725C573,SI1725,end_vn1725);
V1726:VNPU2_2 port map (start_vn,clk,rst,Lc1726,C478V1726,C574V1726,V1726C478,V1726C574,SI1726,end_vn1726);
V1727:VNPU2_2 port map (start_vn,clk,rst,Lc1727,C479V1727,C575V1727,V1727C479,V1727C575,SI1727,end_vn1727);
V1728:VNPU2_2 port map (start_vn,clk,rst,Lc1728,C480V1728,C576V1728,V1728C480,V1728C576,SI1728,end_vn1728);
V1729:VNPU2_2 port map (start_vn,clk,rst,Lc1729,C481V1729,C577V1729,V1729C481,V1729C577,SI1729,end_vn1729);
V1730:VNPU2_2 port map (start_vn,clk,rst,Lc1730,C482V1730,C578V1730,V1730C482,V1730C578,SI1730,end_vn1730);
V1731:VNPU2_2 port map (start_vn,clk,rst,Lc1731,C483V1731,C579V1731,V1731C483,V1731C579,SI1731,end_vn1731);
V1732:VNPU2_2 port map (start_vn,clk,rst,Lc1732,C484V1732,C580V1732,V1732C484,V1732C580,SI1732,end_vn1732);
V1733:VNPU2_2 port map (start_vn,clk,rst,Lc1733,C485V1733,C581V1733,V1733C485,V1733C581,SI1733,end_vn1733);
V1734:VNPU2_2 port map (start_vn,clk,rst,Lc1734,C486V1734,C582V1734,V1734C486,V1734C582,SI1734,end_vn1734);
V1735:VNPU2_2 port map (start_vn,clk,rst,Lc1735,C487V1735,C583V1735,V1735C487,V1735C583,SI1735,end_vn1735);
V1736:VNPU2_2 port map (start_vn,clk,rst,Lc1736,C488V1736,C584V1736,V1736C488,V1736C584,SI1736,end_vn1736);
V1737:VNPU2_2 port map (start_vn,clk,rst,Lc1737,C489V1737,C585V1737,V1737C489,V1737C585,SI1737,end_vn1737);
V1738:VNPU2_2 port map (start_vn,clk,rst,Lc1738,C490V1738,C586V1738,V1738C490,V1738C586,SI1738,end_vn1738);
V1739:VNPU2_2 port map (start_vn,clk,rst,Lc1739,C491V1739,C587V1739,V1739C491,V1739C587,SI1739,end_vn1739);
V1740:VNPU2_2 port map (start_vn,clk,rst,Lc1740,C492V1740,C588V1740,V1740C492,V1740C588,SI1740,end_vn1740);
V1741:VNPU2_2 port map (start_vn,clk,rst,Lc1741,C493V1741,C589V1741,V1741C493,V1741C589,SI1741,end_vn1741);
V1742:VNPU2_2 port map (start_vn,clk,rst,Lc1742,C494V1742,C590V1742,V1742C494,V1742C590,SI1742,end_vn1742);
V1743:VNPU2_2 port map (start_vn,clk,rst,Lc1743,C495V1743,C591V1743,V1743C495,V1743C591,SI1743,end_vn1743);
V1744:VNPU2_2 port map (start_vn,clk,rst,Lc1744,C496V1744,C592V1744,V1744C496,V1744C592,SI1744,end_vn1744);
V1745:VNPU2_2 port map (start_vn,clk,rst,Lc1745,C497V1745,C593V1745,V1745C497,V1745C593,SI1745,end_vn1745);
V1746:VNPU2_2 port map (start_vn,clk,rst,Lc1746,C498V1746,C594V1746,V1746C498,V1746C594,SI1746,end_vn1746);
V1747:VNPU2_2 port map (start_vn,clk,rst,Lc1747,C499V1747,C595V1747,V1747C499,V1747C595,SI1747,end_vn1747);
V1748:VNPU2_2 port map (start_vn,clk,rst,Lc1748,C500V1748,C596V1748,V1748C500,V1748C596,SI1748,end_vn1748);
V1749:VNPU2_2 port map (start_vn,clk,rst,Lc1749,C501V1749,C597V1749,V1749C501,V1749C597,SI1749,end_vn1749);
V1750:VNPU2_2 port map (start_vn,clk,rst,Lc1750,C502V1750,C598V1750,V1750C502,V1750C598,SI1750,end_vn1750);
V1751:VNPU2_2 port map (start_vn,clk,rst,Lc1751,C503V1751,C599V1751,V1751C503,V1751C599,SI1751,end_vn1751);
V1752:VNPU2_2 port map (start_vn,clk,rst,Lc1752,C504V1752,C600V1752,V1752C504,V1752C600,SI1752,end_vn1752);
V1753:VNPU2_2 port map (start_vn,clk,rst,Lc1753,C505V1753,C601V1753,V1753C505,V1753C601,SI1753,end_vn1753);
V1754:VNPU2_2 port map (start_vn,clk,rst,Lc1754,C506V1754,C602V1754,V1754C506,V1754C602,SI1754,end_vn1754);
V1755:VNPU2_2 port map (start_vn,clk,rst,Lc1755,C507V1755,C603V1755,V1755C507,V1755C603,SI1755,end_vn1755);
V1756:VNPU2_2 port map (start_vn,clk,rst,Lc1756,C508V1756,C604V1756,V1756C508,V1756C604,SI1756,end_vn1756);
V1757:VNPU2_2 port map (start_vn,clk,rst,Lc1757,C509V1757,C605V1757,V1757C509,V1757C605,SI1757,end_vn1757);
V1758:VNPU2_2 port map (start_vn,clk,rst,Lc1758,C510V1758,C606V1758,V1758C510,V1758C606,SI1758,end_vn1758);
V1759:VNPU2_2 port map (start_vn,clk,rst,Lc1759,C511V1759,C607V1759,V1759C511,V1759C607,SI1759,end_vn1759);
V1760:VNPU2_2 port map (start_vn,clk,rst,Lc1760,C512V1760,C608V1760,V1760C512,V1760C608,SI1760,end_vn1760);
V1761:VNPU2_2 port map (start_vn,clk,rst,Lc1761,C513V1761,C609V1761,V1761C513,V1761C609,SI1761,end_vn1761);
V1762:VNPU2_2 port map (start_vn,clk,rst,Lc1762,C514V1762,C610V1762,V1762C514,V1762C610,SI1762,end_vn1762);
V1763:VNPU2_2 port map (start_vn,clk,rst,Lc1763,C515V1763,C611V1763,V1763C515,V1763C611,SI1763,end_vn1763);
V1764:VNPU2_2 port map (start_vn,clk,rst,Lc1764,C516V1764,C612V1764,V1764C516,V1764C612,SI1764,end_vn1764);
V1765:VNPU2_2 port map (start_vn,clk,rst,Lc1765,C517V1765,C613V1765,V1765C517,V1765C613,SI1765,end_vn1765);
V1766:VNPU2_2 port map (start_vn,clk,rst,Lc1766,C518V1766,C614V1766,V1766C518,V1766C614,SI1766,end_vn1766);
V1767:VNPU2_2 port map (start_vn,clk,rst,Lc1767,C519V1767,C615V1767,V1767C519,V1767C615,SI1767,end_vn1767);
V1768:VNPU2_2 port map (start_vn,clk,rst,Lc1768,C520V1768,C616V1768,V1768C520,V1768C616,SI1768,end_vn1768);
V1769:VNPU2_2 port map (start_vn,clk,rst,Lc1769,C521V1769,C617V1769,V1769C521,V1769C617,SI1769,end_vn1769);
V1770:VNPU2_2 port map (start_vn,clk,rst,Lc1770,C522V1770,C618V1770,V1770C522,V1770C618,SI1770,end_vn1770);
V1771:VNPU2_2 port map (start_vn,clk,rst,Lc1771,C523V1771,C619V1771,V1771C523,V1771C619,SI1771,end_vn1771);
V1772:VNPU2_2 port map (start_vn,clk,rst,Lc1772,C524V1772,C620V1772,V1772C524,V1772C620,SI1772,end_vn1772);
V1773:VNPU2_2 port map (start_vn,clk,rst,Lc1773,C525V1773,C621V1773,V1773C525,V1773C621,SI1773,end_vn1773);
V1774:VNPU2_2 port map (start_vn,clk,rst,Lc1774,C526V1774,C622V1774,V1774C526,V1774C622,SI1774,end_vn1774);
V1775:VNPU2_2 port map (start_vn,clk,rst,Lc1775,C527V1775,C623V1775,V1775C527,V1775C623,SI1775,end_vn1775);
V1776:VNPU2_2 port map (start_vn,clk,rst,Lc1776,C528V1776,C624V1776,V1776C528,V1776C624,SI1776,end_vn1776);
V1777:VNPU2_2 port map (start_vn,clk,rst,Lc1777,C529V1777,C625V1777,V1777C529,V1777C625,SI1777,end_vn1777);
V1778:VNPU2_2 port map (start_vn,clk,rst,Lc1778,C530V1778,C626V1778,V1778C530,V1778C626,SI1778,end_vn1778);
V1779:VNPU2_2 port map (start_vn,clk,rst,Lc1779,C531V1779,C627V1779,V1779C531,V1779C627,SI1779,end_vn1779);
V1780:VNPU2_2 port map (start_vn,clk,rst,Lc1780,C532V1780,C628V1780,V1780C532,V1780C628,SI1780,end_vn1780);
V1781:VNPU2_2 port map (start_vn,clk,rst,Lc1781,C533V1781,C629V1781,V1781C533,V1781C629,SI1781,end_vn1781);
V1782:VNPU2_2 port map (start_vn,clk,rst,Lc1782,C534V1782,C630V1782,V1782C534,V1782C630,SI1782,end_vn1782);
V1783:VNPU2_2 port map (start_vn,clk,rst,Lc1783,C535V1783,C631V1783,V1783C535,V1783C631,SI1783,end_vn1783);
V1784:VNPU2_2 port map (start_vn,clk,rst,Lc1784,C536V1784,C632V1784,V1784C536,V1784C632,SI1784,end_vn1784);
V1785:VNPU2_2 port map (start_vn,clk,rst,Lc1785,C537V1785,C633V1785,V1785C537,V1785C633,SI1785,end_vn1785);
V1786:VNPU2_2 port map (start_vn,clk,rst,Lc1786,C538V1786,C634V1786,V1786C538,V1786C634,SI1786,end_vn1786);
V1787:VNPU2_2 port map (start_vn,clk,rst,Lc1787,C539V1787,C635V1787,V1787C539,V1787C635,SI1787,end_vn1787);
V1788:VNPU2_2 port map (start_vn,clk,rst,Lc1788,C540V1788,C636V1788,V1788C540,V1788C636,SI1788,end_vn1788);
V1789:VNPU2_2 port map (start_vn,clk,rst,Lc1789,C541V1789,C637V1789,V1789C541,V1789C637,SI1789,end_vn1789);
V1790:VNPU2_2 port map (start_vn,clk,rst,Lc1790,C542V1790,C638V1790,V1790C542,V1790C638,SI1790,end_vn1790);
V1791:VNPU2_2 port map (start_vn,clk,rst,Lc1791,C543V1791,C639V1791,V1791C543,V1791C639,SI1791,end_vn1791);
V1792:VNPU2_2 port map (start_vn,clk,rst,Lc1792,C544V1792,C640V1792,V1792C544,V1792C640,SI1792,end_vn1792);
V1793:VNPU2_2 port map (start_vn,clk,rst,Lc1793,C545V1793,C641V1793,V1793C545,V1793C641,SI1793,end_vn1793);
V1794:VNPU2_2 port map (start_vn,clk,rst,Lc1794,C546V1794,C642V1794,V1794C546,V1794C642,SI1794,end_vn1794);
V1795:VNPU2_2 port map (start_vn,clk,rst,Lc1795,C547V1795,C643V1795,V1795C547,V1795C643,SI1795,end_vn1795);
V1796:VNPU2_2 port map (start_vn,clk,rst,Lc1796,C548V1796,C644V1796,V1796C548,V1796C644,SI1796,end_vn1796);
V1797:VNPU2_2 port map (start_vn,clk,rst,Lc1797,C549V1797,C645V1797,V1797C549,V1797C645,SI1797,end_vn1797);
V1798:VNPU2_2 port map (start_vn,clk,rst,Lc1798,C550V1798,C646V1798,V1798C550,V1798C646,SI1798,end_vn1798);
V1799:VNPU2_2 port map (start_vn,clk,rst,Lc1799,C551V1799,C647V1799,V1799C551,V1799C647,SI1799,end_vn1799);
V1800:VNPU2_2 port map (start_vn,clk,rst,Lc1800,C552V1800,C648V1800,V1800C552,V1800C648,SI1800,end_vn1800);
V1801:VNPU2_2 port map (start_vn,clk,rst,Lc1801,C553V1801,C649V1801,V1801C553,V1801C649,SI1801,end_vn1801);
V1802:VNPU2_2 port map (start_vn,clk,rst,Lc1802,C554V1802,C650V1802,V1802C554,V1802C650,SI1802,end_vn1802);
V1803:VNPU2_2 port map (start_vn,clk,rst,Lc1803,C555V1803,C651V1803,V1803C555,V1803C651,SI1803,end_vn1803);
V1804:VNPU2_2 port map (start_vn,clk,rst,Lc1804,C556V1804,C652V1804,V1804C556,V1804C652,SI1804,end_vn1804);
V1805:VNPU2_2 port map (start_vn,clk,rst,Lc1805,C557V1805,C653V1805,V1805C557,V1805C653,SI1805,end_vn1805);
V1806:VNPU2_2 port map (start_vn,clk,rst,Lc1806,C558V1806,C654V1806,V1806C558,V1806C654,SI1806,end_vn1806);
V1807:VNPU2_2 port map (start_vn,clk,rst,Lc1807,C559V1807,C655V1807,V1807C559,V1807C655,SI1807,end_vn1807);
V1808:VNPU2_2 port map (start_vn,clk,rst,Lc1808,C560V1808,C656V1808,V1808C560,V1808C656,SI1808,end_vn1808);
V1809:VNPU2_2 port map (start_vn,clk,rst,Lc1809,C561V1809,C657V1809,V1809C561,V1809C657,SI1809,end_vn1809);
V1810:VNPU2_2 port map (start_vn,clk,rst,Lc1810,C562V1810,C658V1810,V1810C562,V1810C658,SI1810,end_vn1810);
V1811:VNPU2_2 port map (start_vn,clk,rst,Lc1811,C563V1811,C659V1811,V1811C563,V1811C659,SI1811,end_vn1811);
V1812:VNPU2_2 port map (start_vn,clk,rst,Lc1812,C564V1812,C660V1812,V1812C564,V1812C660,SI1812,end_vn1812);
V1813:VNPU2_2 port map (start_vn,clk,rst,Lc1813,C565V1813,C661V1813,V1813C565,V1813C661,SI1813,end_vn1813);
V1814:VNPU2_2 port map (start_vn,clk,rst,Lc1814,C566V1814,C662V1814,V1814C566,V1814C662,SI1814,end_vn1814);
V1815:VNPU2_2 port map (start_vn,clk,rst,Lc1815,C567V1815,C663V1815,V1815C567,V1815C663,SI1815,end_vn1815);
V1816:VNPU2_2 port map (start_vn,clk,rst,Lc1816,C568V1816,C664V1816,V1816C568,V1816C664,SI1816,end_vn1816);
V1817:VNPU2_2 port map (start_vn,clk,rst,Lc1817,C569V1817,C665V1817,V1817C569,V1817C665,SI1817,end_vn1817);
V1818:VNPU2_2 port map (start_vn,clk,rst,Lc1818,C570V1818,C666V1818,V1818C570,V1818C666,SI1818,end_vn1818);
V1819:VNPU2_2 port map (start_vn,clk,rst,Lc1819,C571V1819,C667V1819,V1819C571,V1819C667,SI1819,end_vn1819);
V1820:VNPU2_2 port map (start_vn,clk,rst,Lc1820,C572V1820,C668V1820,V1820C572,V1820C668,SI1820,end_vn1820);
V1821:VNPU2_2 port map (start_vn,clk,rst,Lc1821,C573V1821,C669V1821,V1821C573,V1821C669,SI1821,end_vn1821);
V1822:VNPU2_2 port map (start_vn,clk,rst,Lc1822,C574V1822,C670V1822,V1822C574,V1822C670,SI1822,end_vn1822);
V1823:VNPU2_2 port map (start_vn,clk,rst,Lc1823,C575V1823,C671V1823,V1823C575,V1823C671,SI1823,end_vn1823);
V1824:VNPU2_2 port map (start_vn,clk,rst,Lc1824,C576V1824,C672V1824,V1824C576,V1824C672,SI1824,end_vn1824);
V1825:VNPU2_2 port map (start_vn,clk,rst,Lc1825,C577V1825,C673V1825,V1825C577,V1825C673,SI1825,end_vn1825);
V1826:VNPU2_2 port map (start_vn,clk,rst,Lc1826,C578V1826,C674V1826,V1826C578,V1826C674,SI1826,end_vn1826);
V1827:VNPU2_2 port map (start_vn,clk,rst,Lc1827,C579V1827,C675V1827,V1827C579,V1827C675,SI1827,end_vn1827);
V1828:VNPU2_2 port map (start_vn,clk,rst,Lc1828,C580V1828,C676V1828,V1828C580,V1828C676,SI1828,end_vn1828);
V1829:VNPU2_2 port map (start_vn,clk,rst,Lc1829,C581V1829,C677V1829,V1829C581,V1829C677,SI1829,end_vn1829);
V1830:VNPU2_2 port map (start_vn,clk,rst,Lc1830,C582V1830,C678V1830,V1830C582,V1830C678,SI1830,end_vn1830);
V1831:VNPU2_2 port map (start_vn,clk,rst,Lc1831,C583V1831,C679V1831,V1831C583,V1831C679,SI1831,end_vn1831);
V1832:VNPU2_2 port map (start_vn,clk,rst,Lc1832,C584V1832,C680V1832,V1832C584,V1832C680,SI1832,end_vn1832);
V1833:VNPU2_2 port map (start_vn,clk,rst,Lc1833,C585V1833,C681V1833,V1833C585,V1833C681,SI1833,end_vn1833);
V1834:VNPU2_2 port map (start_vn,clk,rst,Lc1834,C586V1834,C682V1834,V1834C586,V1834C682,SI1834,end_vn1834);
V1835:VNPU2_2 port map (start_vn,clk,rst,Lc1835,C587V1835,C683V1835,V1835C587,V1835C683,SI1835,end_vn1835);
V1836:VNPU2_2 port map (start_vn,clk,rst,Lc1836,C588V1836,C684V1836,V1836C588,V1836C684,SI1836,end_vn1836);
V1837:VNPU2_2 port map (start_vn,clk,rst,Lc1837,C589V1837,C685V1837,V1837C589,V1837C685,SI1837,end_vn1837);
V1838:VNPU2_2 port map (start_vn,clk,rst,Lc1838,C590V1838,C686V1838,V1838C590,V1838C686,SI1838,end_vn1838);
V1839:VNPU2_2 port map (start_vn,clk,rst,Lc1839,C591V1839,C687V1839,V1839C591,V1839C687,SI1839,end_vn1839);
V1840:VNPU2_2 port map (start_vn,clk,rst,Lc1840,C592V1840,C688V1840,V1840C592,V1840C688,SI1840,end_vn1840);
V1841:VNPU2_2 port map (start_vn,clk,rst,Lc1841,C593V1841,C689V1841,V1841C593,V1841C689,SI1841,end_vn1841);
V1842:VNPU2_2 port map (start_vn,clk,rst,Lc1842,C594V1842,C690V1842,V1842C594,V1842C690,SI1842,end_vn1842);
V1843:VNPU2_2 port map (start_vn,clk,rst,Lc1843,C595V1843,C691V1843,V1843C595,V1843C691,SI1843,end_vn1843);
V1844:VNPU2_2 port map (start_vn,clk,rst,Lc1844,C596V1844,C692V1844,V1844C596,V1844C692,SI1844,end_vn1844);
V1845:VNPU2_2 port map (start_vn,clk,rst,Lc1845,C597V1845,C693V1845,V1845C597,V1845C693,SI1845,end_vn1845);
V1846:VNPU2_2 port map (start_vn,clk,rst,Lc1846,C598V1846,C694V1846,V1846C598,V1846C694,SI1846,end_vn1846);
V1847:VNPU2_2 port map (start_vn,clk,rst,Lc1847,C599V1847,C695V1847,V1847C599,V1847C695,SI1847,end_vn1847);
V1848:VNPU2_2 port map (start_vn,clk,rst,Lc1848,C600V1848,C696V1848,V1848C600,V1848C696,SI1848,end_vn1848);
V1849:VNPU2_2 port map (start_vn,clk,rst,Lc1849,C601V1849,C697V1849,V1849C601,V1849C697,SI1849,end_vn1849);
V1850:VNPU2_2 port map (start_vn,clk,rst,Lc1850,C602V1850,C698V1850,V1850C602,V1850C698,SI1850,end_vn1850);
V1851:VNPU2_2 port map (start_vn,clk,rst,Lc1851,C603V1851,C699V1851,V1851C603,V1851C699,SI1851,end_vn1851);
V1852:VNPU2_2 port map (start_vn,clk,rst,Lc1852,C604V1852,C700V1852,V1852C604,V1852C700,SI1852,end_vn1852);
V1853:VNPU2_2 port map (start_vn,clk,rst,Lc1853,C605V1853,C701V1853,V1853C605,V1853C701,SI1853,end_vn1853);
V1854:VNPU2_2 port map (start_vn,clk,rst,Lc1854,C606V1854,C702V1854,V1854C606,V1854C702,SI1854,end_vn1854);
V1855:VNPU2_2 port map (start_vn,clk,rst,Lc1855,C607V1855,C703V1855,V1855C607,V1855C703,SI1855,end_vn1855);
V1856:VNPU2_2 port map (start_vn,clk,rst,Lc1856,C608V1856,C704V1856,V1856C608,V1856C704,SI1856,end_vn1856);
V1857:VNPU2_2 port map (start_vn,clk,rst,Lc1857,C609V1857,C705V1857,V1857C609,V1857C705,SI1857,end_vn1857);
V1858:VNPU2_2 port map (start_vn,clk,rst,Lc1858,C610V1858,C706V1858,V1858C610,V1858C706,SI1858,end_vn1858);
V1859:VNPU2_2 port map (start_vn,clk,rst,Lc1859,C611V1859,C707V1859,V1859C611,V1859C707,SI1859,end_vn1859);
V1860:VNPU2_2 port map (start_vn,clk,rst,Lc1860,C612V1860,C708V1860,V1860C612,V1860C708,SI1860,end_vn1860);
V1861:VNPU2_2 port map (start_vn,clk,rst,Lc1861,C613V1861,C709V1861,V1861C613,V1861C709,SI1861,end_vn1861);
V1862:VNPU2_2 port map (start_vn,clk,rst,Lc1862,C614V1862,C710V1862,V1862C614,V1862C710,SI1862,end_vn1862);
V1863:VNPU2_2 port map (start_vn,clk,rst,Lc1863,C615V1863,C711V1863,V1863C615,V1863C711,SI1863,end_vn1863);
V1864:VNPU2_2 port map (start_vn,clk,rst,Lc1864,C616V1864,C712V1864,V1864C616,V1864C712,SI1864,end_vn1864);
V1865:VNPU2_2 port map (start_vn,clk,rst,Lc1865,C617V1865,C713V1865,V1865C617,V1865C713,SI1865,end_vn1865);
V1866:VNPU2_2 port map (start_vn,clk,rst,Lc1866,C618V1866,C714V1866,V1866C618,V1866C714,SI1866,end_vn1866);
V1867:VNPU2_2 port map (start_vn,clk,rst,Lc1867,C619V1867,C715V1867,V1867C619,V1867C715,SI1867,end_vn1867);
V1868:VNPU2_2 port map (start_vn,clk,rst,Lc1868,C620V1868,C716V1868,V1868C620,V1868C716,SI1868,end_vn1868);
V1869:VNPU2_2 port map (start_vn,clk,rst,Lc1869,C621V1869,C717V1869,V1869C621,V1869C717,SI1869,end_vn1869);
V1870:VNPU2_2 port map (start_vn,clk,rst,Lc1870,C622V1870,C718V1870,V1870C622,V1870C718,SI1870,end_vn1870);
V1871:VNPU2_2 port map (start_vn,clk,rst,Lc1871,C623V1871,C719V1871,V1871C623,V1871C719,SI1871,end_vn1871);
V1872:VNPU2_2 port map (start_vn,clk,rst,Lc1872,C624V1872,C720V1872,V1872C624,V1872C720,SI1872,end_vn1872);
V1873:VNPU2_2 port map (start_vn,clk,rst,Lc1873,C625V1873,C721V1873,V1873C625,V1873C721,SI1873,end_vn1873);
V1874:VNPU2_2 port map (start_vn,clk,rst,Lc1874,C626V1874,C722V1874,V1874C626,V1874C722,SI1874,end_vn1874);
V1875:VNPU2_2 port map (start_vn,clk,rst,Lc1875,C627V1875,C723V1875,V1875C627,V1875C723,SI1875,end_vn1875);
V1876:VNPU2_2 port map (start_vn,clk,rst,Lc1876,C628V1876,C724V1876,V1876C628,V1876C724,SI1876,end_vn1876);
V1877:VNPU2_2 port map (start_vn,clk,rst,Lc1877,C629V1877,C725V1877,V1877C629,V1877C725,SI1877,end_vn1877);
V1878:VNPU2_2 port map (start_vn,clk,rst,Lc1878,C630V1878,C726V1878,V1878C630,V1878C726,SI1878,end_vn1878);
V1879:VNPU2_2 port map (start_vn,clk,rst,Lc1879,C631V1879,C727V1879,V1879C631,V1879C727,SI1879,end_vn1879);
V1880:VNPU2_2 port map (start_vn,clk,rst,Lc1880,C632V1880,C728V1880,V1880C632,V1880C728,SI1880,end_vn1880);
V1881:VNPU2_2 port map (start_vn,clk,rst,Lc1881,C633V1881,C729V1881,V1881C633,V1881C729,SI1881,end_vn1881);
V1882:VNPU2_2 port map (start_vn,clk,rst,Lc1882,C634V1882,C730V1882,V1882C634,V1882C730,SI1882,end_vn1882);
V1883:VNPU2_2 port map (start_vn,clk,rst,Lc1883,C635V1883,C731V1883,V1883C635,V1883C731,SI1883,end_vn1883);
V1884:VNPU2_2 port map (start_vn,clk,rst,Lc1884,C636V1884,C732V1884,V1884C636,V1884C732,SI1884,end_vn1884);
V1885:VNPU2_2 port map (start_vn,clk,rst,Lc1885,C637V1885,C733V1885,V1885C637,V1885C733,SI1885,end_vn1885);
V1886:VNPU2_2 port map (start_vn,clk,rst,Lc1886,C638V1886,C734V1886,V1886C638,V1886C734,SI1886,end_vn1886);
V1887:VNPU2_2 port map (start_vn,clk,rst,Lc1887,C639V1887,C735V1887,V1887C639,V1887C735,SI1887,end_vn1887);
V1888:VNPU2_2 port map (start_vn,clk,rst,Lc1888,C640V1888,C736V1888,V1888C640,V1888C736,SI1888,end_vn1888);
V1889:VNPU2_2 port map (start_vn,clk,rst,Lc1889,C641V1889,C737V1889,V1889C641,V1889C737,SI1889,end_vn1889);
V1890:VNPU2_2 port map (start_vn,clk,rst,Lc1890,C642V1890,C738V1890,V1890C642,V1890C738,SI1890,end_vn1890);
V1891:VNPU2_2 port map (start_vn,clk,rst,Lc1891,C643V1891,C739V1891,V1891C643,V1891C739,SI1891,end_vn1891);
V1892:VNPU2_2 port map (start_vn,clk,rst,Lc1892,C644V1892,C740V1892,V1892C644,V1892C740,SI1892,end_vn1892);
V1893:VNPU2_2 port map (start_vn,clk,rst,Lc1893,C645V1893,C741V1893,V1893C645,V1893C741,SI1893,end_vn1893);
V1894:VNPU2_2 port map (start_vn,clk,rst,Lc1894,C646V1894,C742V1894,V1894C646,V1894C742,SI1894,end_vn1894);
V1895:VNPU2_2 port map (start_vn,clk,rst,Lc1895,C647V1895,C743V1895,V1895C647,V1895C743,SI1895,end_vn1895);
V1896:VNPU2_2 port map (start_vn,clk,rst,Lc1896,C648V1896,C744V1896,V1896C648,V1896C744,SI1896,end_vn1896);
V1897:VNPU2_2 port map (start_vn,clk,rst,Lc1897,C649V1897,C745V1897,V1897C649,V1897C745,SI1897,end_vn1897);
V1898:VNPU2_2 port map (start_vn,clk,rst,Lc1898,C650V1898,C746V1898,V1898C650,V1898C746,SI1898,end_vn1898);
V1899:VNPU2_2 port map (start_vn,clk,rst,Lc1899,C651V1899,C747V1899,V1899C651,V1899C747,SI1899,end_vn1899);
V1900:VNPU2_2 port map (start_vn,clk,rst,Lc1900,C652V1900,C748V1900,V1900C652,V1900C748,SI1900,end_vn1900);
V1901:VNPU2_2 port map (start_vn,clk,rst,Lc1901,C653V1901,C749V1901,V1901C653,V1901C749,SI1901,end_vn1901);
V1902:VNPU2_2 port map (start_vn,clk,rst,Lc1902,C654V1902,C750V1902,V1902C654,V1902C750,SI1902,end_vn1902);
V1903:VNPU2_2 port map (start_vn,clk,rst,Lc1903,C655V1903,C751V1903,V1903C655,V1903C751,SI1903,end_vn1903);
V1904:VNPU2_2 port map (start_vn,clk,rst,Lc1904,C656V1904,C752V1904,V1904C656,V1904C752,SI1904,end_vn1904);
V1905:VNPU2_2 port map (start_vn,clk,rst,Lc1905,C657V1905,C753V1905,V1905C657,V1905C753,SI1905,end_vn1905);
V1906:VNPU2_2 port map (start_vn,clk,rst,Lc1906,C658V1906,C754V1906,V1906C658,V1906C754,SI1906,end_vn1906);
V1907:VNPU2_2 port map (start_vn,clk,rst,Lc1907,C659V1907,C755V1907,V1907C659,V1907C755,SI1907,end_vn1907);
V1908:VNPU2_2 port map (start_vn,clk,rst,Lc1908,C660V1908,C756V1908,V1908C660,V1908C756,SI1908,end_vn1908);
V1909:VNPU2_2 port map (start_vn,clk,rst,Lc1909,C661V1909,C757V1909,V1909C661,V1909C757,SI1909,end_vn1909);
V1910:VNPU2_2 port map (start_vn,clk,rst,Lc1910,C662V1910,C758V1910,V1910C662,V1910C758,SI1910,end_vn1910);
V1911:VNPU2_2 port map (start_vn,clk,rst,Lc1911,C663V1911,C759V1911,V1911C663,V1911C759,SI1911,end_vn1911);
V1912:VNPU2_2 port map (start_vn,clk,rst,Lc1912,C664V1912,C760V1912,V1912C664,V1912C760,SI1912,end_vn1912);
V1913:VNPU2_2 port map (start_vn,clk,rst,Lc1913,C665V1913,C761V1913,V1913C665,V1913C761,SI1913,end_vn1913);
V1914:VNPU2_2 port map (start_vn,clk,rst,Lc1914,C666V1914,C762V1914,V1914C666,V1914C762,SI1914,end_vn1914);
V1915:VNPU2_2 port map (start_vn,clk,rst,Lc1915,C667V1915,C763V1915,V1915C667,V1915C763,SI1915,end_vn1915);
V1916:VNPU2_2 port map (start_vn,clk,rst,Lc1916,C668V1916,C764V1916,V1916C668,V1916C764,SI1916,end_vn1916);
V1917:VNPU2_2 port map (start_vn,clk,rst,Lc1917,C669V1917,C765V1917,V1917C669,V1917C765,SI1917,end_vn1917);
V1918:VNPU2_2 port map (start_vn,clk,rst,Lc1918,C670V1918,C766V1918,V1918C670,V1918C766,SI1918,end_vn1918);
V1919:VNPU2_2 port map (start_vn,clk,rst,Lc1919,C671V1919,C767V1919,V1919C671,V1919C767,SI1919,end_vn1919);
V1920:VNPU2_2 port map (start_vn,clk,rst,Lc1920,C672V1920,C768V1920,V1920C672,V1920C768,SI1920,end_vn1920);
V1921:VNPU2_2 port map (start_vn,clk,rst,Lc1921,C673V1921,C769V1921,V1921C673,V1921C769,SI1921,end_vn1921);
V1922:VNPU2_2 port map (start_vn,clk,rst,Lc1922,C674V1922,C770V1922,V1922C674,V1922C770,SI1922,end_vn1922);
V1923:VNPU2_2 port map (start_vn,clk,rst,Lc1923,C675V1923,C771V1923,V1923C675,V1923C771,SI1923,end_vn1923);
V1924:VNPU2_2 port map (start_vn,clk,rst,Lc1924,C676V1924,C772V1924,V1924C676,V1924C772,SI1924,end_vn1924);
V1925:VNPU2_2 port map (start_vn,clk,rst,Lc1925,C677V1925,C773V1925,V1925C677,V1925C773,SI1925,end_vn1925);
V1926:VNPU2_2 port map (start_vn,clk,rst,Lc1926,C678V1926,C774V1926,V1926C678,V1926C774,SI1926,end_vn1926);
V1927:VNPU2_2 port map (start_vn,clk,rst,Lc1927,C679V1927,C775V1927,V1927C679,V1927C775,SI1927,end_vn1927);
V1928:VNPU2_2 port map (start_vn,clk,rst,Lc1928,C680V1928,C776V1928,V1928C680,V1928C776,SI1928,end_vn1928);
V1929:VNPU2_2 port map (start_vn,clk,rst,Lc1929,C681V1929,C777V1929,V1929C681,V1929C777,SI1929,end_vn1929);
V1930:VNPU2_2 port map (start_vn,clk,rst,Lc1930,C682V1930,C778V1930,V1930C682,V1930C778,SI1930,end_vn1930);
V1931:VNPU2_2 port map (start_vn,clk,rst,Lc1931,C683V1931,C779V1931,V1931C683,V1931C779,SI1931,end_vn1931);
V1932:VNPU2_2 port map (start_vn,clk,rst,Lc1932,C684V1932,C780V1932,V1932C684,V1932C780,SI1932,end_vn1932);
V1933:VNPU2_2 port map (start_vn,clk,rst,Lc1933,C685V1933,C781V1933,V1933C685,V1933C781,SI1933,end_vn1933);
V1934:VNPU2_2 port map (start_vn,clk,rst,Lc1934,C686V1934,C782V1934,V1934C686,V1934C782,SI1934,end_vn1934);
V1935:VNPU2_2 port map (start_vn,clk,rst,Lc1935,C687V1935,C783V1935,V1935C687,V1935C783,SI1935,end_vn1935);
V1936:VNPU2_2 port map (start_vn,clk,rst,Lc1936,C688V1936,C784V1936,V1936C688,V1936C784,SI1936,end_vn1936);
V1937:VNPU2_2 port map (start_vn,clk,rst,Lc1937,C689V1937,C785V1937,V1937C689,V1937C785,SI1937,end_vn1937);
V1938:VNPU2_2 port map (start_vn,clk,rst,Lc1938,C690V1938,C786V1938,V1938C690,V1938C786,SI1938,end_vn1938);
V1939:VNPU2_2 port map (start_vn,clk,rst,Lc1939,C691V1939,C787V1939,V1939C691,V1939C787,SI1939,end_vn1939);
V1940:VNPU2_2 port map (start_vn,clk,rst,Lc1940,C692V1940,C788V1940,V1940C692,V1940C788,SI1940,end_vn1940);
V1941:VNPU2_2 port map (start_vn,clk,rst,Lc1941,C693V1941,C789V1941,V1941C693,V1941C789,SI1941,end_vn1941);
V1942:VNPU2_2 port map (start_vn,clk,rst,Lc1942,C694V1942,C790V1942,V1942C694,V1942C790,SI1942,end_vn1942);
V1943:VNPU2_2 port map (start_vn,clk,rst,Lc1943,C695V1943,C791V1943,V1943C695,V1943C791,SI1943,end_vn1943);
V1944:VNPU2_2 port map (start_vn,clk,rst,Lc1944,C696V1944,C792V1944,V1944C696,V1944C792,SI1944,end_vn1944);
V1945:VNPU2_2 port map (start_vn,clk,rst,Lc1945,C697V1945,C793V1945,V1945C697,V1945C793,SI1945,end_vn1945);
V1946:VNPU2_2 port map (start_vn,clk,rst,Lc1946,C698V1946,C794V1946,V1946C698,V1946C794,SI1946,end_vn1946);
V1947:VNPU2_2 port map (start_vn,clk,rst,Lc1947,C699V1947,C795V1947,V1947C699,V1947C795,SI1947,end_vn1947);
V1948:VNPU2_2 port map (start_vn,clk,rst,Lc1948,C700V1948,C796V1948,V1948C700,V1948C796,SI1948,end_vn1948);
V1949:VNPU2_2 port map (start_vn,clk,rst,Lc1949,C701V1949,C797V1949,V1949C701,V1949C797,SI1949,end_vn1949);
V1950:VNPU2_2 port map (start_vn,clk,rst,Lc1950,C702V1950,C798V1950,V1950C702,V1950C798,SI1950,end_vn1950);
V1951:VNPU2_2 port map (start_vn,clk,rst,Lc1951,C703V1951,C799V1951,V1951C703,V1951C799,SI1951,end_vn1951);
V1952:VNPU2_2 port map (start_vn,clk,rst,Lc1952,C704V1952,C800V1952,V1952C704,V1952C800,SI1952,end_vn1952);
V1953:VNPU2_2 port map (start_vn,clk,rst,Lc1953,C705V1953,C801V1953,V1953C705,V1953C801,SI1953,end_vn1953);
V1954:VNPU2_2 port map (start_vn,clk,rst,Lc1954,C706V1954,C802V1954,V1954C706,V1954C802,SI1954,end_vn1954);
V1955:VNPU2_2 port map (start_vn,clk,rst,Lc1955,C707V1955,C803V1955,V1955C707,V1955C803,SI1955,end_vn1955);
V1956:VNPU2_2 port map (start_vn,clk,rst,Lc1956,C708V1956,C804V1956,V1956C708,V1956C804,SI1956,end_vn1956);
V1957:VNPU2_2 port map (start_vn,clk,rst,Lc1957,C709V1957,C805V1957,V1957C709,V1957C805,SI1957,end_vn1957);
V1958:VNPU2_2 port map (start_vn,clk,rst,Lc1958,C710V1958,C806V1958,V1958C710,V1958C806,SI1958,end_vn1958);
V1959:VNPU2_2 port map (start_vn,clk,rst,Lc1959,C711V1959,C807V1959,V1959C711,V1959C807,SI1959,end_vn1959);
V1960:VNPU2_2 port map (start_vn,clk,rst,Lc1960,C712V1960,C808V1960,V1960C712,V1960C808,SI1960,end_vn1960);
V1961:VNPU2_2 port map (start_vn,clk,rst,Lc1961,C713V1961,C809V1961,V1961C713,V1961C809,SI1961,end_vn1961);
V1962:VNPU2_2 port map (start_vn,clk,rst,Lc1962,C714V1962,C810V1962,V1962C714,V1962C810,SI1962,end_vn1962);
V1963:VNPU2_2 port map (start_vn,clk,rst,Lc1963,C715V1963,C811V1963,V1963C715,V1963C811,SI1963,end_vn1963);
V1964:VNPU2_2 port map (start_vn,clk,rst,Lc1964,C716V1964,C812V1964,V1964C716,V1964C812,SI1964,end_vn1964);
V1965:VNPU2_2 port map (start_vn,clk,rst,Lc1965,C717V1965,C813V1965,V1965C717,V1965C813,SI1965,end_vn1965);
V1966:VNPU2_2 port map (start_vn,clk,rst,Lc1966,C718V1966,C814V1966,V1966C718,V1966C814,SI1966,end_vn1966);
V1967:VNPU2_2 port map (start_vn,clk,rst,Lc1967,C719V1967,C815V1967,V1967C719,V1967C815,SI1967,end_vn1967);
V1968:VNPU2_2 port map (start_vn,clk,rst,Lc1968,C720V1968,C816V1968,V1968C720,V1968C816,SI1968,end_vn1968);
V1969:VNPU2_2 port map (start_vn,clk,rst,Lc1969,C721V1969,C817V1969,V1969C721,V1969C817,SI1969,end_vn1969);
V1970:VNPU2_2 port map (start_vn,clk,rst,Lc1970,C722V1970,C818V1970,V1970C722,V1970C818,SI1970,end_vn1970);
V1971:VNPU2_2 port map (start_vn,clk,rst,Lc1971,C723V1971,C819V1971,V1971C723,V1971C819,SI1971,end_vn1971);
V1972:VNPU2_2 port map (start_vn,clk,rst,Lc1972,C724V1972,C820V1972,V1972C724,V1972C820,SI1972,end_vn1972);
V1973:VNPU2_2 port map (start_vn,clk,rst,Lc1973,C725V1973,C821V1973,V1973C725,V1973C821,SI1973,end_vn1973);
V1974:VNPU2_2 port map (start_vn,clk,rst,Lc1974,C726V1974,C822V1974,V1974C726,V1974C822,SI1974,end_vn1974);
V1975:VNPU2_2 port map (start_vn,clk,rst,Lc1975,C727V1975,C823V1975,V1975C727,V1975C823,SI1975,end_vn1975);
V1976:VNPU2_2 port map (start_vn,clk,rst,Lc1976,C728V1976,C824V1976,V1976C728,V1976C824,SI1976,end_vn1976);
V1977:VNPU2_2 port map (start_vn,clk,rst,Lc1977,C729V1977,C825V1977,V1977C729,V1977C825,SI1977,end_vn1977);
V1978:VNPU2_2 port map (start_vn,clk,rst,Lc1978,C730V1978,C826V1978,V1978C730,V1978C826,SI1978,end_vn1978);
V1979:VNPU2_2 port map (start_vn,clk,rst,Lc1979,C731V1979,C827V1979,V1979C731,V1979C827,SI1979,end_vn1979);
V1980:VNPU2_2 port map (start_vn,clk,rst,Lc1980,C732V1980,C828V1980,V1980C732,V1980C828,SI1980,end_vn1980);
V1981:VNPU2_2 port map (start_vn,clk,rst,Lc1981,C733V1981,C829V1981,V1981C733,V1981C829,SI1981,end_vn1981);
V1982:VNPU2_2 port map (start_vn,clk,rst,Lc1982,C734V1982,C830V1982,V1982C734,V1982C830,SI1982,end_vn1982);
V1983:VNPU2_2 port map (start_vn,clk,rst,Lc1983,C735V1983,C831V1983,V1983C735,V1983C831,SI1983,end_vn1983);
V1984:VNPU2_2 port map (start_vn,clk,rst,Lc1984,C736V1984,C832V1984,V1984C736,V1984C832,SI1984,end_vn1984);
V1985:VNPU2_2 port map (start_vn,clk,rst,Lc1985,C737V1985,C833V1985,V1985C737,V1985C833,SI1985,end_vn1985);
V1986:VNPU2_2 port map (start_vn,clk,rst,Lc1986,C738V1986,C834V1986,V1986C738,V1986C834,SI1986,end_vn1986);
V1987:VNPU2_2 port map (start_vn,clk,rst,Lc1987,C739V1987,C835V1987,V1987C739,V1987C835,SI1987,end_vn1987);
V1988:VNPU2_2 port map (start_vn,clk,rst,Lc1988,C740V1988,C836V1988,V1988C740,V1988C836,SI1988,end_vn1988);
V1989:VNPU2_2 port map (start_vn,clk,rst,Lc1989,C741V1989,C837V1989,V1989C741,V1989C837,SI1989,end_vn1989);
V1990:VNPU2_2 port map (start_vn,clk,rst,Lc1990,C742V1990,C838V1990,V1990C742,V1990C838,SI1990,end_vn1990);
V1991:VNPU2_2 port map (start_vn,clk,rst,Lc1991,C743V1991,C839V1991,V1991C743,V1991C839,SI1991,end_vn1991);
V1992:VNPU2_2 port map (start_vn,clk,rst,Lc1992,C744V1992,C840V1992,V1992C744,V1992C840,SI1992,end_vn1992);
V1993:VNPU2_2 port map (start_vn,clk,rst,Lc1993,C745V1993,C841V1993,V1993C745,V1993C841,SI1993,end_vn1993);
V1994:VNPU2_2 port map (start_vn,clk,rst,Lc1994,C746V1994,C842V1994,V1994C746,V1994C842,SI1994,end_vn1994);
V1995:VNPU2_2 port map (start_vn,clk,rst,Lc1995,C747V1995,C843V1995,V1995C747,V1995C843,SI1995,end_vn1995);
V1996:VNPU2_2 port map (start_vn,clk,rst,Lc1996,C748V1996,C844V1996,V1996C748,V1996C844,SI1996,end_vn1996);
V1997:VNPU2_2 port map (start_vn,clk,rst,Lc1997,C749V1997,C845V1997,V1997C749,V1997C845,SI1997,end_vn1997);
V1998:VNPU2_2 port map (start_vn,clk,rst,Lc1998,C750V1998,C846V1998,V1998C750,V1998C846,SI1998,end_vn1998);
V1999:VNPU2_2 port map (start_vn,clk,rst,Lc1999,C751V1999,C847V1999,V1999C751,V1999C847,SI1999,end_vn1999);
V2000:VNPU2_2 port map (start_vn,clk,rst,Lc2000,C752V2000,C848V2000,V2000C752,V2000C848,SI2000,end_vn2000);
V2001:VNPU2_2 port map (start_vn,clk,rst,Lc2001,C753V2001,C849V2001,V2001C753,V2001C849,SI2001,end_vn2001);
V2002:VNPU2_2 port map (start_vn,clk,rst,Lc2002,C754V2002,C850V2002,V2002C754,V2002C850,SI2002,end_vn2002);
V2003:VNPU2_2 port map (start_vn,clk,rst,Lc2003,C755V2003,C851V2003,V2003C755,V2003C851,SI2003,end_vn2003);
V2004:VNPU2_2 port map (start_vn,clk,rst,Lc2004,C756V2004,C852V2004,V2004C756,V2004C852,SI2004,end_vn2004);
V2005:VNPU2_2 port map (start_vn,clk,rst,Lc2005,C757V2005,C853V2005,V2005C757,V2005C853,SI2005,end_vn2005);
V2006:VNPU2_2 port map (start_vn,clk,rst,Lc2006,C758V2006,C854V2006,V2006C758,V2006C854,SI2006,end_vn2006);
V2007:VNPU2_2 port map (start_vn,clk,rst,Lc2007,C759V2007,C855V2007,V2007C759,V2007C855,SI2007,end_vn2007);
V2008:VNPU2_2 port map (start_vn,clk,rst,Lc2008,C760V2008,C856V2008,V2008C760,V2008C856,SI2008,end_vn2008);
V2009:VNPU2_2 port map (start_vn,clk,rst,Lc2009,C761V2009,C857V2009,V2009C761,V2009C857,SI2009,end_vn2009);
V2010:VNPU2_2 port map (start_vn,clk,rst,Lc2010,C762V2010,C858V2010,V2010C762,V2010C858,SI2010,end_vn2010);
V2011:VNPU2_2 port map (start_vn,clk,rst,Lc2011,C763V2011,C859V2011,V2011C763,V2011C859,SI2011,end_vn2011);
V2012:VNPU2_2 port map (start_vn,clk,rst,Lc2012,C764V2012,C860V2012,V2012C764,V2012C860,SI2012,end_vn2012);
V2013:VNPU2_2 port map (start_vn,clk,rst,Lc2013,C765V2013,C861V2013,V2013C765,V2013C861,SI2013,end_vn2013);
V2014:VNPU2_2 port map (start_vn,clk,rst,Lc2014,C766V2014,C862V2014,V2014C766,V2014C862,SI2014,end_vn2014);
V2015:VNPU2_2 port map (start_vn,clk,rst,Lc2015,C767V2015,C863V2015,V2015C767,V2015C863,SI2015,end_vn2015);
V2016:VNPU2_2 port map (start_vn,clk,rst,Lc2016,C768V2016,C864V2016,V2016C768,V2016C864,SI2016,end_vn2016);
V2017:VNPU2_2 port map (start_vn,clk,rst,Lc2017,C769V2017,C865V2017,V2017C769,V2017C865,SI2017,end_vn2017);
V2018:VNPU2_2 port map (start_vn,clk,rst,Lc2018,C770V2018,C866V2018,V2018C770,V2018C866,SI2018,end_vn2018);
V2019:VNPU2_2 port map (start_vn,clk,rst,Lc2019,C771V2019,C867V2019,V2019C771,V2019C867,SI2019,end_vn2019);
V2020:VNPU2_2 port map (start_vn,clk,rst,Lc2020,C772V2020,C868V2020,V2020C772,V2020C868,SI2020,end_vn2020);
V2021:VNPU2_2 port map (start_vn,clk,rst,Lc2021,C773V2021,C869V2021,V2021C773,V2021C869,SI2021,end_vn2021);
V2022:VNPU2_2 port map (start_vn,clk,rst,Lc2022,C774V2022,C870V2022,V2022C774,V2022C870,SI2022,end_vn2022);
V2023:VNPU2_2 port map (start_vn,clk,rst,Lc2023,C775V2023,C871V2023,V2023C775,V2023C871,SI2023,end_vn2023);
V2024:VNPU2_2 port map (start_vn,clk,rst,Lc2024,C776V2024,C872V2024,V2024C776,V2024C872,SI2024,end_vn2024);
V2025:VNPU2_2 port map (start_vn,clk,rst,Lc2025,C777V2025,C873V2025,V2025C777,V2025C873,SI2025,end_vn2025);
V2026:VNPU2_2 port map (start_vn,clk,rst,Lc2026,C778V2026,C874V2026,V2026C778,V2026C874,SI2026,end_vn2026);
V2027:VNPU2_2 port map (start_vn,clk,rst,Lc2027,C779V2027,C875V2027,V2027C779,V2027C875,SI2027,end_vn2027);
V2028:VNPU2_2 port map (start_vn,clk,rst,Lc2028,C780V2028,C876V2028,V2028C780,V2028C876,SI2028,end_vn2028);
V2029:VNPU2_2 port map (start_vn,clk,rst,Lc2029,C781V2029,C877V2029,V2029C781,V2029C877,SI2029,end_vn2029);
V2030:VNPU2_2 port map (start_vn,clk,rst,Lc2030,C782V2030,C878V2030,V2030C782,V2030C878,SI2030,end_vn2030);
V2031:VNPU2_2 port map (start_vn,clk,rst,Lc2031,C783V2031,C879V2031,V2031C783,V2031C879,SI2031,end_vn2031);
V2032:VNPU2_2 port map (start_vn,clk,rst,Lc2032,C784V2032,C880V2032,V2032C784,V2032C880,SI2032,end_vn2032);
V2033:VNPU2_2 port map (start_vn,clk,rst,Lc2033,C785V2033,C881V2033,V2033C785,V2033C881,SI2033,end_vn2033);
V2034:VNPU2_2 port map (start_vn,clk,rst,Lc2034,C786V2034,C882V2034,V2034C786,V2034C882,SI2034,end_vn2034);
V2035:VNPU2_2 port map (start_vn,clk,rst,Lc2035,C787V2035,C883V2035,V2035C787,V2035C883,SI2035,end_vn2035);
V2036:VNPU2_2 port map (start_vn,clk,rst,Lc2036,C788V2036,C884V2036,V2036C788,V2036C884,SI2036,end_vn2036);
V2037:VNPU2_2 port map (start_vn,clk,rst,Lc2037,C789V2037,C885V2037,V2037C789,V2037C885,SI2037,end_vn2037);
V2038:VNPU2_2 port map (start_vn,clk,rst,Lc2038,C790V2038,C886V2038,V2038C790,V2038C886,SI2038,end_vn2038);
V2039:VNPU2_2 port map (start_vn,clk,rst,Lc2039,C791V2039,C887V2039,V2039C791,V2039C887,SI2039,end_vn2039);
V2040:VNPU2_2 port map (start_vn,clk,rst,Lc2040,C792V2040,C888V2040,V2040C792,V2040C888,SI2040,end_vn2040);
V2041:VNPU2_2 port map (start_vn,clk,rst,Lc2041,C793V2041,C889V2041,V2041C793,V2041C889,SI2041,end_vn2041);
V2042:VNPU2_2 port map (start_vn,clk,rst,Lc2042,C794V2042,C890V2042,V2042C794,V2042C890,SI2042,end_vn2042);
V2043:VNPU2_2 port map (start_vn,clk,rst,Lc2043,C795V2043,C891V2043,V2043C795,V2043C891,SI2043,end_vn2043);
V2044:VNPU2_2 port map (start_vn,clk,rst,Lc2044,C796V2044,C892V2044,V2044C796,V2044C892,SI2044,end_vn2044);
V2045:VNPU2_2 port map (start_vn,clk,rst,Lc2045,C797V2045,C893V2045,V2045C797,V2045C893,SI2045,end_vn2045);
V2046:VNPU2_2 port map (start_vn,clk,rst,Lc2046,C798V2046,C894V2046,V2046C798,V2046C894,SI2046,end_vn2046);
V2047:VNPU2_2 port map (start_vn,clk,rst,Lc2047,C799V2047,C895V2047,V2047C799,V2047C895,SI2047,end_vn2047);
V2048:VNPU2_2 port map (start_vn,clk,rst,Lc2048,C800V2048,C896V2048,V2048C800,V2048C896,SI2048,end_vn2048);
V2049:VNPU2_2 port map (start_vn,clk,rst,Lc2049,C801V2049,C897V2049,V2049C801,V2049C897,SI2049,end_vn2049);
V2050:VNPU2_2 port map (start_vn,clk,rst,Lc2050,C802V2050,C898V2050,V2050C802,V2050C898,SI2050,end_vn2050);
V2051:VNPU2_2 port map (start_vn,clk,rst,Lc2051,C803V2051,C899V2051,V2051C803,V2051C899,SI2051,end_vn2051);
V2052:VNPU2_2 port map (start_vn,clk,rst,Lc2052,C804V2052,C900V2052,V2052C804,V2052C900,SI2052,end_vn2052);
V2053:VNPU2_2 port map (start_vn,clk,rst,Lc2053,C805V2053,C901V2053,V2053C805,V2053C901,SI2053,end_vn2053);
V2054:VNPU2_2 port map (start_vn,clk,rst,Lc2054,C806V2054,C902V2054,V2054C806,V2054C902,SI2054,end_vn2054);
V2055:VNPU2_2 port map (start_vn,clk,rst,Lc2055,C807V2055,C903V2055,V2055C807,V2055C903,SI2055,end_vn2055);
V2056:VNPU2_2 port map (start_vn,clk,rst,Lc2056,C808V2056,C904V2056,V2056C808,V2056C904,SI2056,end_vn2056);
V2057:VNPU2_2 port map (start_vn,clk,rst,Lc2057,C809V2057,C905V2057,V2057C809,V2057C905,SI2057,end_vn2057);
V2058:VNPU2_2 port map (start_vn,clk,rst,Lc2058,C810V2058,C906V2058,V2058C810,V2058C906,SI2058,end_vn2058);
V2059:VNPU2_2 port map (start_vn,clk,rst,Lc2059,C811V2059,C907V2059,V2059C811,V2059C907,SI2059,end_vn2059);
V2060:VNPU2_2 port map (start_vn,clk,rst,Lc2060,C812V2060,C908V2060,V2060C812,V2060C908,SI2060,end_vn2060);
V2061:VNPU2_2 port map (start_vn,clk,rst,Lc2061,C813V2061,C909V2061,V2061C813,V2061C909,SI2061,end_vn2061);
V2062:VNPU2_2 port map (start_vn,clk,rst,Lc2062,C814V2062,C910V2062,V2062C814,V2062C910,SI2062,end_vn2062);
V2063:VNPU2_2 port map (start_vn,clk,rst,Lc2063,C815V2063,C911V2063,V2063C815,V2063C911,SI2063,end_vn2063);
V2064:VNPU2_2 port map (start_vn,clk,rst,Lc2064,C816V2064,C912V2064,V2064C816,V2064C912,SI2064,end_vn2064);
V2065:VNPU2_2 port map (start_vn,clk,rst,Lc2065,C817V2065,C913V2065,V2065C817,V2065C913,SI2065,end_vn2065);
V2066:VNPU2_2 port map (start_vn,clk,rst,Lc2066,C818V2066,C914V2066,V2066C818,V2066C914,SI2066,end_vn2066);
V2067:VNPU2_2 port map (start_vn,clk,rst,Lc2067,C819V2067,C915V2067,V2067C819,V2067C915,SI2067,end_vn2067);
V2068:VNPU2_2 port map (start_vn,clk,rst,Lc2068,C820V2068,C916V2068,V2068C820,V2068C916,SI2068,end_vn2068);
V2069:VNPU2_2 port map (start_vn,clk,rst,Lc2069,C821V2069,C917V2069,V2069C821,V2069C917,SI2069,end_vn2069);
V2070:VNPU2_2 port map (start_vn,clk,rst,Lc2070,C822V2070,C918V2070,V2070C822,V2070C918,SI2070,end_vn2070);
V2071:VNPU2_2 port map (start_vn,clk,rst,Lc2071,C823V2071,C919V2071,V2071C823,V2071C919,SI2071,end_vn2071);
V2072:VNPU2_2 port map (start_vn,clk,rst,Lc2072,C824V2072,C920V2072,V2072C824,V2072C920,SI2072,end_vn2072);
V2073:VNPU2_2 port map (start_vn,clk,rst,Lc2073,C825V2073,C921V2073,V2073C825,V2073C921,SI2073,end_vn2073);
V2074:VNPU2_2 port map (start_vn,clk,rst,Lc2074,C826V2074,C922V2074,V2074C826,V2074C922,SI2074,end_vn2074);
V2075:VNPU2_2 port map (start_vn,clk,rst,Lc2075,C827V2075,C923V2075,V2075C827,V2075C923,SI2075,end_vn2075);
V2076:VNPU2_2 port map (start_vn,clk,rst,Lc2076,C828V2076,C924V2076,V2076C828,V2076C924,SI2076,end_vn2076);
V2077:VNPU2_2 port map (start_vn,clk,rst,Lc2077,C829V2077,C925V2077,V2077C829,V2077C925,SI2077,end_vn2077);
V2078:VNPU2_2 port map (start_vn,clk,rst,Lc2078,C830V2078,C926V2078,V2078C830,V2078C926,SI2078,end_vn2078);
V2079:VNPU2_2 port map (start_vn,clk,rst,Lc2079,C831V2079,C927V2079,V2079C831,V2079C927,SI2079,end_vn2079);
V2080:VNPU2_2 port map (start_vn,clk,rst,Lc2080,C832V2080,C928V2080,V2080C832,V2080C928,SI2080,end_vn2080);
V2081:VNPU2_2 port map (start_vn,clk,rst,Lc2081,C833V2081,C929V2081,V2081C833,V2081C929,SI2081,end_vn2081);
V2082:VNPU2_2 port map (start_vn,clk,rst,Lc2082,C834V2082,C930V2082,V2082C834,V2082C930,SI2082,end_vn2082);
V2083:VNPU2_2 port map (start_vn,clk,rst,Lc2083,C835V2083,C931V2083,V2083C835,V2083C931,SI2083,end_vn2083);
V2084:VNPU2_2 port map (start_vn,clk,rst,Lc2084,C836V2084,C932V2084,V2084C836,V2084C932,SI2084,end_vn2084);
V2085:VNPU2_2 port map (start_vn,clk,rst,Lc2085,C837V2085,C933V2085,V2085C837,V2085C933,SI2085,end_vn2085);
V2086:VNPU2_2 port map (start_vn,clk,rst,Lc2086,C838V2086,C934V2086,V2086C838,V2086C934,SI2086,end_vn2086);
V2087:VNPU2_2 port map (start_vn,clk,rst,Lc2087,C839V2087,C935V2087,V2087C839,V2087C935,SI2087,end_vn2087);
V2088:VNPU2_2 port map (start_vn,clk,rst,Lc2088,C840V2088,C936V2088,V2088C840,V2088C936,SI2088,end_vn2088);
V2089:VNPU2_2 port map (start_vn,clk,rst,Lc2089,C841V2089,C937V2089,V2089C841,V2089C937,SI2089,end_vn2089);
V2090:VNPU2_2 port map (start_vn,clk,rst,Lc2090,C842V2090,C938V2090,V2090C842,V2090C938,SI2090,end_vn2090);
V2091:VNPU2_2 port map (start_vn,clk,rst,Lc2091,C843V2091,C939V2091,V2091C843,V2091C939,SI2091,end_vn2091);
V2092:VNPU2_2 port map (start_vn,clk,rst,Lc2092,C844V2092,C940V2092,V2092C844,V2092C940,SI2092,end_vn2092);
V2093:VNPU2_2 port map (start_vn,clk,rst,Lc2093,C845V2093,C941V2093,V2093C845,V2093C941,SI2093,end_vn2093);
V2094:VNPU2_2 port map (start_vn,clk,rst,Lc2094,C846V2094,C942V2094,V2094C846,V2094C942,SI2094,end_vn2094);
V2095:VNPU2_2 port map (start_vn,clk,rst,Lc2095,C847V2095,C943V2095,V2095C847,V2095C943,SI2095,end_vn2095);
V2096:VNPU2_2 port map (start_vn,clk,rst,Lc2096,C848V2096,C944V2096,V2096C848,V2096C944,SI2096,end_vn2096);
V2097:VNPU2_2 port map (start_vn,clk,rst,Lc2097,C849V2097,C945V2097,V2097C849,V2097C945,SI2097,end_vn2097);
V2098:VNPU2_2 port map (start_vn,clk,rst,Lc2098,C850V2098,C946V2098,V2098C850,V2098C946,SI2098,end_vn2098);
V2099:VNPU2_2 port map (start_vn,clk,rst,Lc2099,C851V2099,C947V2099,V2099C851,V2099C947,SI2099,end_vn2099);
V2100:VNPU2_2 port map (start_vn,clk,rst,Lc2100,C852V2100,C948V2100,V2100C852,V2100C948,SI2100,end_vn2100);
V2101:VNPU2_2 port map (start_vn,clk,rst,Lc2101,C853V2101,C949V2101,V2101C853,V2101C949,SI2101,end_vn2101);
V2102:VNPU2_2 port map (start_vn,clk,rst,Lc2102,C854V2102,C950V2102,V2102C854,V2102C950,SI2102,end_vn2102);
V2103:VNPU2_2 port map (start_vn,clk,rst,Lc2103,C855V2103,C951V2103,V2103C855,V2103C951,SI2103,end_vn2103);
V2104:VNPU2_2 port map (start_vn,clk,rst,Lc2104,C856V2104,C952V2104,V2104C856,V2104C952,SI2104,end_vn2104);
V2105:VNPU2_2 port map (start_vn,clk,rst,Lc2105,C857V2105,C953V2105,V2105C857,V2105C953,SI2105,end_vn2105);
V2106:VNPU2_2 port map (start_vn,clk,rst,Lc2106,C858V2106,C954V2106,V2106C858,V2106C954,SI2106,end_vn2106);
V2107:VNPU2_2 port map (start_vn,clk,rst,Lc2107,C859V2107,C955V2107,V2107C859,V2107C955,SI2107,end_vn2107);
V2108:VNPU2_2 port map (start_vn,clk,rst,Lc2108,C860V2108,C956V2108,V2108C860,V2108C956,SI2108,end_vn2108);
V2109:VNPU2_2 port map (start_vn,clk,rst,Lc2109,C861V2109,C957V2109,V2109C861,V2109C957,SI2109,end_vn2109);
V2110:VNPU2_2 port map (start_vn,clk,rst,Lc2110,C862V2110,C958V2110,V2110C862,V2110C958,SI2110,end_vn2110);
V2111:VNPU2_2 port map (start_vn,clk,rst,Lc2111,C863V2111,C959V2111,V2111C863,V2111C959,SI2111,end_vn2111);
V2112:VNPU2_2 port map (start_vn,clk,rst,Lc2112,C864V2112,C960V2112,V2112C864,V2112C960,SI2112,end_vn2112);
V2113:VNPU2_2 port map (start_vn,clk,rst,Lc2113,C865V2113,C961V2113,V2113C865,V2113C961,SI2113,end_vn2113);
V2114:VNPU2_2 port map (start_vn,clk,rst,Lc2114,C866V2114,C962V2114,V2114C866,V2114C962,SI2114,end_vn2114);
V2115:VNPU2_2 port map (start_vn,clk,rst,Lc2115,C867V2115,C963V2115,V2115C867,V2115C963,SI2115,end_vn2115);
V2116:VNPU2_2 port map (start_vn,clk,rst,Lc2116,C868V2116,C964V2116,V2116C868,V2116C964,SI2116,end_vn2116);
V2117:VNPU2_2 port map (start_vn,clk,rst,Lc2117,C869V2117,C965V2117,V2117C869,V2117C965,SI2117,end_vn2117);
V2118:VNPU2_2 port map (start_vn,clk,rst,Lc2118,C870V2118,C966V2118,V2118C870,V2118C966,SI2118,end_vn2118);
V2119:VNPU2_2 port map (start_vn,clk,rst,Lc2119,C871V2119,C967V2119,V2119C871,V2119C967,SI2119,end_vn2119);
V2120:VNPU2_2 port map (start_vn,clk,rst,Lc2120,C872V2120,C968V2120,V2120C872,V2120C968,SI2120,end_vn2120);
V2121:VNPU2_2 port map (start_vn,clk,rst,Lc2121,C873V2121,C969V2121,V2121C873,V2121C969,SI2121,end_vn2121);
V2122:VNPU2_2 port map (start_vn,clk,rst,Lc2122,C874V2122,C970V2122,V2122C874,V2122C970,SI2122,end_vn2122);
V2123:VNPU2_2 port map (start_vn,clk,rst,Lc2123,C875V2123,C971V2123,V2123C875,V2123C971,SI2123,end_vn2123);
V2124:VNPU2_2 port map (start_vn,clk,rst,Lc2124,C876V2124,C972V2124,V2124C876,V2124C972,SI2124,end_vn2124);
V2125:VNPU2_2 port map (start_vn,clk,rst,Lc2125,C877V2125,C973V2125,V2125C877,V2125C973,SI2125,end_vn2125);
V2126:VNPU2_2 port map (start_vn,clk,rst,Lc2126,C878V2126,C974V2126,V2126C878,V2126C974,SI2126,end_vn2126);
V2127:VNPU2_2 port map (start_vn,clk,rst,Lc2127,C879V2127,C975V2127,V2127C879,V2127C975,SI2127,end_vn2127);
V2128:VNPU2_2 port map (start_vn,clk,rst,Lc2128,C880V2128,C976V2128,V2128C880,V2128C976,SI2128,end_vn2128);
V2129:VNPU2_2 port map (start_vn,clk,rst,Lc2129,C881V2129,C977V2129,V2129C881,V2129C977,SI2129,end_vn2129);
V2130:VNPU2_2 port map (start_vn,clk,rst,Lc2130,C882V2130,C978V2130,V2130C882,V2130C978,SI2130,end_vn2130);
V2131:VNPU2_2 port map (start_vn,clk,rst,Lc2131,C883V2131,C979V2131,V2131C883,V2131C979,SI2131,end_vn2131);
V2132:VNPU2_2 port map (start_vn,clk,rst,Lc2132,C884V2132,C980V2132,V2132C884,V2132C980,SI2132,end_vn2132);
V2133:VNPU2_2 port map (start_vn,clk,rst,Lc2133,C885V2133,C981V2133,V2133C885,V2133C981,SI2133,end_vn2133);
V2134:VNPU2_2 port map (start_vn,clk,rst,Lc2134,C886V2134,C982V2134,V2134C886,V2134C982,SI2134,end_vn2134);
V2135:VNPU2_2 port map (start_vn,clk,rst,Lc2135,C887V2135,C983V2135,V2135C887,V2135C983,SI2135,end_vn2135);
V2136:VNPU2_2 port map (start_vn,clk,rst,Lc2136,C888V2136,C984V2136,V2136C888,V2136C984,SI2136,end_vn2136);
V2137:VNPU2_2 port map (start_vn,clk,rst,Lc2137,C889V2137,C985V2137,V2137C889,V2137C985,SI2137,end_vn2137);
V2138:VNPU2_2 port map (start_vn,clk,rst,Lc2138,C890V2138,C986V2138,V2138C890,V2138C986,SI2138,end_vn2138);
V2139:VNPU2_2 port map (start_vn,clk,rst,Lc2139,C891V2139,C987V2139,V2139C891,V2139C987,SI2139,end_vn2139);
V2140:VNPU2_2 port map (start_vn,clk,rst,Lc2140,C892V2140,C988V2140,V2140C892,V2140C988,SI2140,end_vn2140);
V2141:VNPU2_2 port map (start_vn,clk,rst,Lc2141,C893V2141,C989V2141,V2141C893,V2141C989,SI2141,end_vn2141);
V2142:VNPU2_2 port map (start_vn,clk,rst,Lc2142,C894V2142,C990V2142,V2142C894,V2142C990,SI2142,end_vn2142);
V2143:VNPU2_2 port map (start_vn,clk,rst,Lc2143,C895V2143,C991V2143,V2143C895,V2143C991,SI2143,end_vn2143);
V2144:VNPU2_2 port map (start_vn,clk,rst,Lc2144,C896V2144,C992V2144,V2144C896,V2144C992,SI2144,end_vn2144);
V2145:VNPU2_2 port map (start_vn,clk,rst,Lc2145,C897V2145,C993V2145,V2145C897,V2145C993,SI2145,end_vn2145);
V2146:VNPU2_2 port map (start_vn,clk,rst,Lc2146,C898V2146,C994V2146,V2146C898,V2146C994,SI2146,end_vn2146);
V2147:VNPU2_2 port map (start_vn,clk,rst,Lc2147,C899V2147,C995V2147,V2147C899,V2147C995,SI2147,end_vn2147);
V2148:VNPU2_2 port map (start_vn,clk,rst,Lc2148,C900V2148,C996V2148,V2148C900,V2148C996,SI2148,end_vn2148);
V2149:VNPU2_2 port map (start_vn,clk,rst,Lc2149,C901V2149,C997V2149,V2149C901,V2149C997,SI2149,end_vn2149);
V2150:VNPU2_2 port map (start_vn,clk,rst,Lc2150,C902V2150,C998V2150,V2150C902,V2150C998,SI2150,end_vn2150);
V2151:VNPU2_2 port map (start_vn,clk,rst,Lc2151,C903V2151,C999V2151,V2151C903,V2151C999,SI2151,end_vn2151);
V2152:VNPU2_2 port map (start_vn,clk,rst,Lc2152,C904V2152,C1000V2152,V2152C904,V2152C1000,SI2152,end_vn2152);
V2153:VNPU2_2 port map (start_vn,clk,rst,Lc2153,C905V2153,C1001V2153,V2153C905,V2153C1001,SI2153,end_vn2153);
V2154:VNPU2_2 port map (start_vn,clk,rst,Lc2154,C906V2154,C1002V2154,V2154C906,V2154C1002,SI2154,end_vn2154);
V2155:VNPU2_2 port map (start_vn,clk,rst,Lc2155,C907V2155,C1003V2155,V2155C907,V2155C1003,SI2155,end_vn2155);
V2156:VNPU2_2 port map (start_vn,clk,rst,Lc2156,C908V2156,C1004V2156,V2156C908,V2156C1004,SI2156,end_vn2156);
V2157:VNPU2_2 port map (start_vn,clk,rst,Lc2157,C909V2157,C1005V2157,V2157C909,V2157C1005,SI2157,end_vn2157);
V2158:VNPU2_2 port map (start_vn,clk,rst,Lc2158,C910V2158,C1006V2158,V2158C910,V2158C1006,SI2158,end_vn2158);
V2159:VNPU2_2 port map (start_vn,clk,rst,Lc2159,C911V2159,C1007V2159,V2159C911,V2159C1007,SI2159,end_vn2159);
V2160:VNPU2_2 port map (start_vn,clk,rst,Lc2160,C912V2160,C1008V2160,V2160C912,V2160C1008,SI2160,end_vn2160);
V2161:VNPU2_2 port map (start_vn,clk,rst,Lc2161,C913V2161,C1009V2161,V2161C913,V2161C1009,SI2161,end_vn2161);
V2162:VNPU2_2 port map (start_vn,clk,rst,Lc2162,C914V2162,C1010V2162,V2162C914,V2162C1010,SI2162,end_vn2162);
V2163:VNPU2_2 port map (start_vn,clk,rst,Lc2163,C915V2163,C1011V2163,V2163C915,V2163C1011,SI2163,end_vn2163);
V2164:VNPU2_2 port map (start_vn,clk,rst,Lc2164,C916V2164,C1012V2164,V2164C916,V2164C1012,SI2164,end_vn2164);
V2165:VNPU2_2 port map (start_vn,clk,rst,Lc2165,C917V2165,C1013V2165,V2165C917,V2165C1013,SI2165,end_vn2165);
V2166:VNPU2_2 port map (start_vn,clk,rst,Lc2166,C918V2166,C1014V2166,V2166C918,V2166C1014,SI2166,end_vn2166);
V2167:VNPU2_2 port map (start_vn,clk,rst,Lc2167,C919V2167,C1015V2167,V2167C919,V2167C1015,SI2167,end_vn2167);
V2168:VNPU2_2 port map (start_vn,clk,rst,Lc2168,C920V2168,C1016V2168,V2168C920,V2168C1016,SI2168,end_vn2168);
V2169:VNPU2_2 port map (start_vn,clk,rst,Lc2169,C921V2169,C1017V2169,V2169C921,V2169C1017,SI2169,end_vn2169);
V2170:VNPU2_2 port map (start_vn,clk,rst,Lc2170,C922V2170,C1018V2170,V2170C922,V2170C1018,SI2170,end_vn2170);
V2171:VNPU2_2 port map (start_vn,clk,rst,Lc2171,C923V2171,C1019V2171,V2171C923,V2171C1019,SI2171,end_vn2171);
V2172:VNPU2_2 port map (start_vn,clk,rst,Lc2172,C924V2172,C1020V2172,V2172C924,V2172C1020,SI2172,end_vn2172);
V2173:VNPU2_2 port map (start_vn,clk,rst,Lc2173,C925V2173,C1021V2173,V2173C925,V2173C1021,SI2173,end_vn2173);
V2174:VNPU2_2 port map (start_vn,clk,rst,Lc2174,C926V2174,C1022V2174,V2174C926,V2174C1022,SI2174,end_vn2174);
V2175:VNPU2_2 port map (start_vn,clk,rst,Lc2175,C927V2175,C1023V2175,V2175C927,V2175C1023,SI2175,end_vn2175);
V2176:VNPU2_2 port map (start_vn,clk,rst,Lc2176,C928V2176,C1024V2176,V2176C928,V2176C1024,SI2176,end_vn2176);
V2177:VNPU2_2 port map (start_vn,clk,rst,Lc2177,C929V2177,C1025V2177,V2177C929,V2177C1025,SI2177,end_vn2177);
V2178:VNPU2_2 port map (start_vn,clk,rst,Lc2178,C930V2178,C1026V2178,V2178C930,V2178C1026,SI2178,end_vn2178);
V2179:VNPU2_2 port map (start_vn,clk,rst,Lc2179,C931V2179,C1027V2179,V2179C931,V2179C1027,SI2179,end_vn2179);
V2180:VNPU2_2 port map (start_vn,clk,rst,Lc2180,C932V2180,C1028V2180,V2180C932,V2180C1028,SI2180,end_vn2180);
V2181:VNPU2_2 port map (start_vn,clk,rst,Lc2181,C933V2181,C1029V2181,V2181C933,V2181C1029,SI2181,end_vn2181);
V2182:VNPU2_2 port map (start_vn,clk,rst,Lc2182,C934V2182,C1030V2182,V2182C934,V2182C1030,SI2182,end_vn2182);
V2183:VNPU2_2 port map (start_vn,clk,rst,Lc2183,C935V2183,C1031V2183,V2183C935,V2183C1031,SI2183,end_vn2183);
V2184:VNPU2_2 port map (start_vn,clk,rst,Lc2184,C936V2184,C1032V2184,V2184C936,V2184C1032,SI2184,end_vn2184);
V2185:VNPU2_2 port map (start_vn,clk,rst,Lc2185,C937V2185,C1033V2185,V2185C937,V2185C1033,SI2185,end_vn2185);
V2186:VNPU2_2 port map (start_vn,clk,rst,Lc2186,C938V2186,C1034V2186,V2186C938,V2186C1034,SI2186,end_vn2186);
V2187:VNPU2_2 port map (start_vn,clk,rst,Lc2187,C939V2187,C1035V2187,V2187C939,V2187C1035,SI2187,end_vn2187);
V2188:VNPU2_2 port map (start_vn,clk,rst,Lc2188,C940V2188,C1036V2188,V2188C940,V2188C1036,SI2188,end_vn2188);
V2189:VNPU2_2 port map (start_vn,clk,rst,Lc2189,C941V2189,C1037V2189,V2189C941,V2189C1037,SI2189,end_vn2189);
V2190:VNPU2_2 port map (start_vn,clk,rst,Lc2190,C942V2190,C1038V2190,V2190C942,V2190C1038,SI2190,end_vn2190);
V2191:VNPU2_2 port map (start_vn,clk,rst,Lc2191,C943V2191,C1039V2191,V2191C943,V2191C1039,SI2191,end_vn2191);
V2192:VNPU2_2 port map (start_vn,clk,rst,Lc2192,C944V2192,C1040V2192,V2192C944,V2192C1040,SI2192,end_vn2192);
V2193:VNPU2_2 port map (start_vn,clk,rst,Lc2193,C945V2193,C1041V2193,V2193C945,V2193C1041,SI2193,end_vn2193);
V2194:VNPU2_2 port map (start_vn,clk,rst,Lc2194,C946V2194,C1042V2194,V2194C946,V2194C1042,SI2194,end_vn2194);
V2195:VNPU2_2 port map (start_vn,clk,rst,Lc2195,C947V2195,C1043V2195,V2195C947,V2195C1043,SI2195,end_vn2195);
V2196:VNPU2_2 port map (start_vn,clk,rst,Lc2196,C948V2196,C1044V2196,V2196C948,V2196C1044,SI2196,end_vn2196);
V2197:VNPU2_2 port map (start_vn,clk,rst,Lc2197,C949V2197,C1045V2197,V2197C949,V2197C1045,SI2197,end_vn2197);
V2198:VNPU2_2 port map (start_vn,clk,rst,Lc2198,C950V2198,C1046V2198,V2198C950,V2198C1046,SI2198,end_vn2198);
V2199:VNPU2_2 port map (start_vn,clk,rst,Lc2199,C951V2199,C1047V2199,V2199C951,V2199C1047,SI2199,end_vn2199);
V2200:VNPU2_2 port map (start_vn,clk,rst,Lc2200,C952V2200,C1048V2200,V2200C952,V2200C1048,SI2200,end_vn2200);
V2201:VNPU2_2 port map (start_vn,clk,rst,Lc2201,C953V2201,C1049V2201,V2201C953,V2201C1049,SI2201,end_vn2201);
V2202:VNPU2_2 port map (start_vn,clk,rst,Lc2202,C954V2202,C1050V2202,V2202C954,V2202C1050,SI2202,end_vn2202);
V2203:VNPU2_2 port map (start_vn,clk,rst,Lc2203,C955V2203,C1051V2203,V2203C955,V2203C1051,SI2203,end_vn2203);
V2204:VNPU2_2 port map (start_vn,clk,rst,Lc2204,C956V2204,C1052V2204,V2204C956,V2204C1052,SI2204,end_vn2204);
V2205:VNPU2_2 port map (start_vn,clk,rst,Lc2205,C957V2205,C1053V2205,V2205C957,V2205C1053,SI2205,end_vn2205);
V2206:VNPU2_2 port map (start_vn,clk,rst,Lc2206,C958V2206,C1054V2206,V2206C958,V2206C1054,SI2206,end_vn2206);
V2207:VNPU2_2 port map (start_vn,clk,rst,Lc2207,C959V2207,C1055V2207,V2207C959,V2207C1055,SI2207,end_vn2207);
V2208:VNPU2_2 port map (start_vn,clk,rst,Lc2208,C960V2208,C1056V2208,V2208C960,V2208C1056,SI2208,end_vn2208);
V2209:VNPU2_2 port map (start_vn,clk,rst,Lc2209,C961V2209,C1057V2209,V2209C961,V2209C1057,SI2209,end_vn2209);
V2210:VNPU2_2 port map (start_vn,clk,rst,Lc2210,C962V2210,C1058V2210,V2210C962,V2210C1058,SI2210,end_vn2210);
V2211:VNPU2_2 port map (start_vn,clk,rst,Lc2211,C963V2211,C1059V2211,V2211C963,V2211C1059,SI2211,end_vn2211);
V2212:VNPU2_2 port map (start_vn,clk,rst,Lc2212,C964V2212,C1060V2212,V2212C964,V2212C1060,SI2212,end_vn2212);
V2213:VNPU2_2 port map (start_vn,clk,rst,Lc2213,C965V2213,C1061V2213,V2213C965,V2213C1061,SI2213,end_vn2213);
V2214:VNPU2_2 port map (start_vn,clk,rst,Lc2214,C966V2214,C1062V2214,V2214C966,V2214C1062,SI2214,end_vn2214);
V2215:VNPU2_2 port map (start_vn,clk,rst,Lc2215,C967V2215,C1063V2215,V2215C967,V2215C1063,SI2215,end_vn2215);
V2216:VNPU2_2 port map (start_vn,clk,rst,Lc2216,C968V2216,C1064V2216,V2216C968,V2216C1064,SI2216,end_vn2216);
V2217:VNPU2_2 port map (start_vn,clk,rst,Lc2217,C969V2217,C1065V2217,V2217C969,V2217C1065,SI2217,end_vn2217);
V2218:VNPU2_2 port map (start_vn,clk,rst,Lc2218,C970V2218,C1066V2218,V2218C970,V2218C1066,SI2218,end_vn2218);
V2219:VNPU2_2 port map (start_vn,clk,rst,Lc2219,C971V2219,C1067V2219,V2219C971,V2219C1067,SI2219,end_vn2219);
V2220:VNPU2_2 port map (start_vn,clk,rst,Lc2220,C972V2220,C1068V2220,V2220C972,V2220C1068,SI2220,end_vn2220);
V2221:VNPU2_2 port map (start_vn,clk,rst,Lc2221,C973V2221,C1069V2221,V2221C973,V2221C1069,SI2221,end_vn2221);
V2222:VNPU2_2 port map (start_vn,clk,rst,Lc2222,C974V2222,C1070V2222,V2222C974,V2222C1070,SI2222,end_vn2222);
V2223:VNPU2_2 port map (start_vn,clk,rst,Lc2223,C975V2223,C1071V2223,V2223C975,V2223C1071,SI2223,end_vn2223);
V2224:VNPU2_2 port map (start_vn,clk,rst,Lc2224,C976V2224,C1072V2224,V2224C976,V2224C1072,SI2224,end_vn2224);
V2225:VNPU2_2 port map (start_vn,clk,rst,Lc2225,C977V2225,C1073V2225,V2225C977,V2225C1073,SI2225,end_vn2225);
V2226:VNPU2_2 port map (start_vn,clk,rst,Lc2226,C978V2226,C1074V2226,V2226C978,V2226C1074,SI2226,end_vn2226);
V2227:VNPU2_2 port map (start_vn,clk,rst,Lc2227,C979V2227,C1075V2227,V2227C979,V2227C1075,SI2227,end_vn2227);
V2228:VNPU2_2 port map (start_vn,clk,rst,Lc2228,C980V2228,C1076V2228,V2228C980,V2228C1076,SI2228,end_vn2228);
V2229:VNPU2_2 port map (start_vn,clk,rst,Lc2229,C981V2229,C1077V2229,V2229C981,V2229C1077,SI2229,end_vn2229);
V2230:VNPU2_2 port map (start_vn,clk,rst,Lc2230,C982V2230,C1078V2230,V2230C982,V2230C1078,SI2230,end_vn2230);
V2231:VNPU2_2 port map (start_vn,clk,rst,Lc2231,C983V2231,C1079V2231,V2231C983,V2231C1079,SI2231,end_vn2231);
V2232:VNPU2_2 port map (start_vn,clk,rst,Lc2232,C984V2232,C1080V2232,V2232C984,V2232C1080,SI2232,end_vn2232);
V2233:VNPU2_2 port map (start_vn,clk,rst,Lc2233,C985V2233,C1081V2233,V2233C985,V2233C1081,SI2233,end_vn2233);
V2234:VNPU2_2 port map (start_vn,clk,rst,Lc2234,C986V2234,C1082V2234,V2234C986,V2234C1082,SI2234,end_vn2234);
V2235:VNPU2_2 port map (start_vn,clk,rst,Lc2235,C987V2235,C1083V2235,V2235C987,V2235C1083,SI2235,end_vn2235);
V2236:VNPU2_2 port map (start_vn,clk,rst,Lc2236,C988V2236,C1084V2236,V2236C988,V2236C1084,SI2236,end_vn2236);
V2237:VNPU2_2 port map (start_vn,clk,rst,Lc2237,C989V2237,C1085V2237,V2237C989,V2237C1085,SI2237,end_vn2237);
V2238:VNPU2_2 port map (start_vn,clk,rst,Lc2238,C990V2238,C1086V2238,V2238C990,V2238C1086,SI2238,end_vn2238);
V2239:VNPU2_2 port map (start_vn,clk,rst,Lc2239,C991V2239,C1087V2239,V2239C991,V2239C1087,SI2239,end_vn2239);
V2240:VNPU2_2 port map (start_vn,clk,rst,Lc2240,C992V2240,C1088V2240,V2240C992,V2240C1088,SI2240,end_vn2240);
V2241:VNPU2_2 port map (start_vn,clk,rst,Lc2241,C993V2241,C1089V2241,V2241C993,V2241C1089,SI2241,end_vn2241);
V2242:VNPU2_2 port map (start_vn,clk,rst,Lc2242,C994V2242,C1090V2242,V2242C994,V2242C1090,SI2242,end_vn2242);
V2243:VNPU2_2 port map (start_vn,clk,rst,Lc2243,C995V2243,C1091V2243,V2243C995,V2243C1091,SI2243,end_vn2243);
V2244:VNPU2_2 port map (start_vn,clk,rst,Lc2244,C996V2244,C1092V2244,V2244C996,V2244C1092,SI2244,end_vn2244);
V2245:VNPU2_2 port map (start_vn,clk,rst,Lc2245,C997V2245,C1093V2245,V2245C997,V2245C1093,SI2245,end_vn2245);
V2246:VNPU2_2 port map (start_vn,clk,rst,Lc2246,C998V2246,C1094V2246,V2246C998,V2246C1094,SI2246,end_vn2246);
V2247:VNPU2_2 port map (start_vn,clk,rst,Lc2247,C999V2247,C1095V2247,V2247C999,V2247C1095,SI2247,end_vn2247);
V2248:VNPU2_2 port map (start_vn,clk,rst,Lc2248,C1000V2248,C1096V2248,V2248C1000,V2248C1096,SI2248,end_vn2248);
V2249:VNPU2_2 port map (start_vn,clk,rst,Lc2249,C1001V2249,C1097V2249,V2249C1001,V2249C1097,SI2249,end_vn2249);
V2250:VNPU2_2 port map (start_vn,clk,rst,Lc2250,C1002V2250,C1098V2250,V2250C1002,V2250C1098,SI2250,end_vn2250);
V2251:VNPU2_2 port map (start_vn,clk,rst,Lc2251,C1003V2251,C1099V2251,V2251C1003,V2251C1099,SI2251,end_vn2251);
V2252:VNPU2_2 port map (start_vn,clk,rst,Lc2252,C1004V2252,C1100V2252,V2252C1004,V2252C1100,SI2252,end_vn2252);
V2253:VNPU2_2 port map (start_vn,clk,rst,Lc2253,C1005V2253,C1101V2253,V2253C1005,V2253C1101,SI2253,end_vn2253);
V2254:VNPU2_2 port map (start_vn,clk,rst,Lc2254,C1006V2254,C1102V2254,V2254C1006,V2254C1102,SI2254,end_vn2254);
V2255:VNPU2_2 port map (start_vn,clk,rst,Lc2255,C1007V2255,C1103V2255,V2255C1007,V2255C1103,SI2255,end_vn2255);
V2256:VNPU2_2 port map (start_vn,clk,rst,Lc2256,C1008V2256,C1104V2256,V2256C1008,V2256C1104,SI2256,end_vn2256);
V2257:VNPU2_2 port map (start_vn,clk,rst,Lc2257,C1009V2257,C1105V2257,V2257C1009,V2257C1105,SI2257,end_vn2257);
V2258:VNPU2_2 port map (start_vn,clk,rst,Lc2258,C1010V2258,C1106V2258,V2258C1010,V2258C1106,SI2258,end_vn2258);
V2259:VNPU2_2 port map (start_vn,clk,rst,Lc2259,C1011V2259,C1107V2259,V2259C1011,V2259C1107,SI2259,end_vn2259);
V2260:VNPU2_2 port map (start_vn,clk,rst,Lc2260,C1012V2260,C1108V2260,V2260C1012,V2260C1108,SI2260,end_vn2260);
V2261:VNPU2_2 port map (start_vn,clk,rst,Lc2261,C1013V2261,C1109V2261,V2261C1013,V2261C1109,SI2261,end_vn2261);
V2262:VNPU2_2 port map (start_vn,clk,rst,Lc2262,C1014V2262,C1110V2262,V2262C1014,V2262C1110,SI2262,end_vn2262);
V2263:VNPU2_2 port map (start_vn,clk,rst,Lc2263,C1015V2263,C1111V2263,V2263C1015,V2263C1111,SI2263,end_vn2263);
V2264:VNPU2_2 port map (start_vn,clk,rst,Lc2264,C1016V2264,C1112V2264,V2264C1016,V2264C1112,SI2264,end_vn2264);
V2265:VNPU2_2 port map (start_vn,clk,rst,Lc2265,C1017V2265,C1113V2265,V2265C1017,V2265C1113,SI2265,end_vn2265);
V2266:VNPU2_2 port map (start_vn,clk,rst,Lc2266,C1018V2266,C1114V2266,V2266C1018,V2266C1114,SI2266,end_vn2266);
V2267:VNPU2_2 port map (start_vn,clk,rst,Lc2267,C1019V2267,C1115V2267,V2267C1019,V2267C1115,SI2267,end_vn2267);
V2268:VNPU2_2 port map (start_vn,clk,rst,Lc2268,C1020V2268,C1116V2268,V2268C1020,V2268C1116,SI2268,end_vn2268);
V2269:VNPU2_2 port map (start_vn,clk,rst,Lc2269,C1021V2269,C1117V2269,V2269C1021,V2269C1117,SI2269,end_vn2269);
V2270:VNPU2_2 port map (start_vn,clk,rst,Lc2270,C1022V2270,C1118V2270,V2270C1022,V2270C1118,SI2270,end_vn2270);
V2271:VNPU2_2 port map (start_vn,clk,rst,Lc2271,C1023V2271,C1119V2271,V2271C1023,V2271C1119,SI2271,end_vn2271);
V2272:VNPU2_2 port map (start_vn,clk,rst,Lc2272,C1024V2272,C1120V2272,V2272C1024,V2272C1120,SI2272,end_vn2272);
V2273:VNPU2_2 port map (start_vn,clk,rst,Lc2273,C1025V2273,C1121V2273,V2273C1025,V2273C1121,SI2273,end_vn2273);
V2274:VNPU2_2 port map (start_vn,clk,rst,Lc2274,C1026V2274,C1122V2274,V2274C1026,V2274C1122,SI2274,end_vn2274);
V2275:VNPU2_2 port map (start_vn,clk,rst,Lc2275,C1027V2275,C1123V2275,V2275C1027,V2275C1123,SI2275,end_vn2275);
V2276:VNPU2_2 port map (start_vn,clk,rst,Lc2276,C1028V2276,C1124V2276,V2276C1028,V2276C1124,SI2276,end_vn2276);
V2277:VNPU2_2 port map (start_vn,clk,rst,Lc2277,C1029V2277,C1125V2277,V2277C1029,V2277C1125,SI2277,end_vn2277);
V2278:VNPU2_2 port map (start_vn,clk,rst,Lc2278,C1030V2278,C1126V2278,V2278C1030,V2278C1126,SI2278,end_vn2278);
V2279:VNPU2_2 port map (start_vn,clk,rst,Lc2279,C1031V2279,C1127V2279,V2279C1031,V2279C1127,SI2279,end_vn2279);
V2280:VNPU2_2 port map (start_vn,clk,rst,Lc2280,C1032V2280,C1128V2280,V2280C1032,V2280C1128,SI2280,end_vn2280);
V2281:VNPU2_2 port map (start_vn,clk,rst,Lc2281,C1033V2281,C1129V2281,V2281C1033,V2281C1129,SI2281,end_vn2281);
V2282:VNPU2_2 port map (start_vn,clk,rst,Lc2282,C1034V2282,C1130V2282,V2282C1034,V2282C1130,SI2282,end_vn2282);
V2283:VNPU2_2 port map (start_vn,clk,rst,Lc2283,C1035V2283,C1131V2283,V2283C1035,V2283C1131,SI2283,end_vn2283);
V2284:VNPU2_2 port map (start_vn,clk,rst,Lc2284,C1036V2284,C1132V2284,V2284C1036,V2284C1132,SI2284,end_vn2284);
V2285:VNPU2_2 port map (start_vn,clk,rst,Lc2285,C1037V2285,C1133V2285,V2285C1037,V2285C1133,SI2285,end_vn2285);
V2286:VNPU2_2 port map (start_vn,clk,rst,Lc2286,C1038V2286,C1134V2286,V2286C1038,V2286C1134,SI2286,end_vn2286);
V2287:VNPU2_2 port map (start_vn,clk,rst,Lc2287,C1039V2287,C1135V2287,V2287C1039,V2287C1135,SI2287,end_vn2287);
V2288:VNPU2_2 port map (start_vn,clk,rst,Lc2288,C1040V2288,C1136V2288,V2288C1040,V2288C1136,SI2288,end_vn2288);
V2289:VNPU2_2 port map (start_vn,clk,rst,Lc2289,C1041V2289,C1137V2289,V2289C1041,V2289C1137,SI2289,end_vn2289);
V2290:VNPU2_2 port map (start_vn,clk,rst,Lc2290,C1042V2290,C1138V2290,V2290C1042,V2290C1138,SI2290,end_vn2290);
V2291:VNPU2_2 port map (start_vn,clk,rst,Lc2291,C1043V2291,C1139V2291,V2291C1043,V2291C1139,SI2291,end_vn2291);
V2292:VNPU2_2 port map (start_vn,clk,rst,Lc2292,C1044V2292,C1140V2292,V2292C1044,V2292C1140,SI2292,end_vn2292);
V2293:VNPU2_2 port map (start_vn,clk,rst,Lc2293,C1045V2293,C1141V2293,V2293C1045,V2293C1141,SI2293,end_vn2293);
V2294:VNPU2_2 port map (start_vn,clk,rst,Lc2294,C1046V2294,C1142V2294,V2294C1046,V2294C1142,SI2294,end_vn2294);
V2295:VNPU2_2 port map (start_vn,clk,rst,Lc2295,C1047V2295,C1143V2295,V2295C1047,V2295C1143,SI2295,end_vn2295);
V2296:VNPU2_2 port map (start_vn,clk,rst,Lc2296,C1048V2296,C1144V2296,V2296C1048,V2296C1144,SI2296,end_vn2296);
V2297:VNPU2_2 port map (start_vn,clk,rst,Lc2297,C1049V2297,C1145V2297,V2297C1049,V2297C1145,SI2297,end_vn2297);
V2298:VNPU2_2 port map (start_vn,clk,rst,Lc2298,C1050V2298,C1146V2298,V2298C1050,V2298C1146,SI2298,end_vn2298);
V2299:VNPU2_2 port map (start_vn,clk,rst,Lc2299,C1051V2299,C1147V2299,V2299C1051,V2299C1147,SI2299,end_vn2299);
V2300:VNPU2_2 port map (start_vn,clk,rst,Lc2300,C1052V2300,C1148V2300,V2300C1052,V2300C1148,SI2300,end_vn2300);
V2301:VNPU2_2 port map (start_vn,clk,rst,Lc2301,C1053V2301,C1149V2301,V2301C1053,V2301C1149,SI2301,end_vn2301);
V2302:VNPU2_2 port map (start_vn,clk,rst,Lc2302,C1054V2302,C1150V2302,V2302C1054,V2302C1150,SI2302,end_vn2302);
V2303:VNPU2_2 port map (start_vn,clk,rst,Lc2303,C1055V2303,C1151V2303,V2303C1055,V2303C1151,SI2303,end_vn2303);
V2304:VNPU2_2 port map (start_vn,clk,rst,Lc2304,C1056V2304,C1152V2304,V2304C1056,V2304C1152,SI2304,end_vn2304);
end_cnt<=end_cn1 and end_cn2 and end_cn3 and end_cn4 and end_cn5 and end_cn6 and end_cn7 and end_cn8 and end_cn9 and end_cn10 and end_cn11 and end_cn12 and end_cn13 and end_cn14 and end_cn15 and end_cn16 and end_cn17 and end_cn18 and end_cn19 and end_cn20 and end_cn21 and end_cn22 and end_cn23 and end_cn24 and end_cn25 and end_cn26 and end_cn27 and end_cn28 and end_cn29 and end_cn30 and end_cn31 and end_cn32 and end_cn33 and end_cn34 and end_cn35 and end_cn36 and end_cn37 and end_cn38 and end_cn39 and end_cn40 and end_cn41 and end_cn42 and end_cn43 and end_cn44 and end_cn45 and end_cn46 and end_cn47 and end_cn48 and end_cn49 and end_cn50 and end_cn51 and end_cn52 and end_cn53 and end_cn54 and end_cn55 and end_cn56 and end_cn57 and end_cn58 and end_cn59 and end_cn60 and end_cn61 and end_cn62 and end_cn63 and end_cn64 and end_cn65 and end_cn66 and end_cn67 and end_cn68 and end_cn69 and end_cn70 and end_cn71 and end_cn72 and end_cn73 and end_cn74 and end_cn75 and end_cn76 and end_cn77 and end_cn78 and end_cn79 and end_cn80 and end_cn81 and end_cn82 and end_cn83 and end_cn84 and end_cn85 and end_cn86 and end_cn87 and end_cn88 and end_cn89 and end_cn90 and end_cn91 and end_cn92 and end_cn93 and end_cn94 and end_cn95 and end_cn96 and end_cn97 and end_cn98 and end_cn99 and end_cn100 and end_cn101 and end_cn102 and end_cn103 and end_cn104 and end_cn105 and end_cn106 and end_cn107 and end_cn108 and end_cn109 and end_cn110 and end_cn111 and end_cn112 and end_cn113 and end_cn114 and end_cn115 and end_cn116 and end_cn117 and end_cn118 and end_cn119 and end_cn120 and end_cn121 and end_cn122 and end_cn123 and end_cn124 and end_cn125 and end_cn126 and end_cn127 and end_cn128 and end_cn129 and end_cn130 and end_cn131 and end_cn132 and end_cn133 and end_cn134 and end_cn135 and end_cn136 and end_cn137 and end_cn138 and end_cn139 and end_cn140 and end_cn141 and end_cn142 and end_cn143 and end_cn144 and end_cn145 and end_cn146 and end_cn147 and end_cn148 and end_cn149 and end_cn150 and end_cn151 and end_cn152 and end_cn153 and end_cn154 and end_cn155 and end_cn156 and end_cn157 and end_cn158 and end_cn159 and end_cn160 and end_cn161 and end_cn162 and end_cn163 and end_cn164 and end_cn165 and end_cn166 and end_cn167 and end_cn168 and end_cn169 and end_cn170 and end_cn171 and end_cn172 and end_cn173 and end_cn174 and end_cn175 and end_cn176 and end_cn177 and end_cn178 and end_cn179 and end_cn180 and end_cn181 and end_cn182 and end_cn183 and end_cn184 and end_cn185 and end_cn186 and end_cn187 and end_cn188 and end_cn189 and end_cn190 and end_cn191 and end_cn192 and end_cn193 and end_cn194 and end_cn195 and end_cn196 and end_cn197 and end_cn198 and end_cn199 and end_cn200 and end_cn201 and end_cn202 and end_cn203 and end_cn204 and end_cn205 and end_cn206 and end_cn207 and end_cn208 and end_cn209 and end_cn210 and end_cn211 and end_cn212 and end_cn213 and end_cn214 and end_cn215 and end_cn216 and end_cn217 and end_cn218 and end_cn219 and end_cn220 and end_cn221 and end_cn222 and end_cn223 and end_cn224 and end_cn225 and end_cn226 and end_cn227 and end_cn228 and end_cn229 and end_cn230 and end_cn231 and end_cn232 and end_cn233 and end_cn234 and end_cn235 and end_cn236 and end_cn237 and end_cn238 and end_cn239 and end_cn240 and end_cn241 and end_cn242 and end_cn243 and end_cn244 and end_cn245 and end_cn246 and end_cn247 and end_cn248 and end_cn249 and end_cn250 and end_cn251 and end_cn252 and end_cn253 and end_cn254 and end_cn255 and end_cn256 and end_cn257 and end_cn258 and end_cn259 and end_cn260 and end_cn261 and end_cn262 and end_cn263 and end_cn264 and end_cn265 and end_cn266 and end_cn267 and end_cn268 and end_cn269 and end_cn270 and end_cn271 and end_cn272 and end_cn273 and end_cn274 and end_cn275 and end_cn276 and end_cn277 and end_cn278 and end_cn279 and end_cn280 and end_cn281 and end_cn282 and end_cn283 and end_cn284 and end_cn285 and end_cn286 and end_cn287 and end_cn288 and end_cn289 and end_cn290 and end_cn291 and end_cn292 and end_cn293 and end_cn294 and end_cn295 and end_cn296 and end_cn297 and end_cn298 and end_cn299 and end_cn300 and end_cn301 and end_cn302 and end_cn303 and end_cn304 and end_cn305 and end_cn306 and end_cn307 and end_cn308 and end_cn309 and end_cn310 and end_cn311 and end_cn312 and end_cn313 and end_cn314 and end_cn315 and end_cn316 and end_cn317 and end_cn318 and end_cn319 and end_cn320 and end_cn321 and end_cn322 and end_cn323 and end_cn324 and end_cn325 and end_cn326 and end_cn327 and end_cn328 and end_cn329 and end_cn330 and end_cn331 and end_cn332 and end_cn333 and end_cn334 and end_cn335 and end_cn336 and end_cn337 and end_cn338 and end_cn339 and end_cn340 and end_cn341 and end_cn342 and end_cn343 and end_cn344 and end_cn345 and end_cn346 and end_cn347 and end_cn348 and end_cn349 and end_cn350 and end_cn351 and end_cn352 and end_cn353 and end_cn354 and end_cn355 and end_cn356 and end_cn357 and end_cn358 and end_cn359 and end_cn360 and end_cn361 and end_cn362 and end_cn363 and end_cn364 and end_cn365 and end_cn366 and end_cn367 and end_cn368 and end_cn369 and end_cn370 and end_cn371 and end_cn372 and end_cn373 and end_cn374 and end_cn375 and end_cn376 and end_cn377 and end_cn378 and end_cn379 and end_cn380 and end_cn381 and end_cn382 and end_cn383 and end_cn384 and end_cn385 and end_cn386 and end_cn387 and end_cn388 and end_cn389 and end_cn390 and end_cn391 and end_cn392 and end_cn393 and end_cn394 and end_cn395 and end_cn396 and end_cn397 and end_cn398 and end_cn399 and end_cn400 and end_cn401 and end_cn402 and end_cn403 and end_cn404 and end_cn405 and end_cn406 and end_cn407 and end_cn408 and end_cn409 and end_cn410 and end_cn411 and end_cn412 and end_cn413 and end_cn414 and end_cn415 and end_cn416 and end_cn417 and end_cn418 and end_cn419 and end_cn420 and end_cn421 and end_cn422 and end_cn423 and end_cn424 and end_cn425 and end_cn426 and end_cn427 and end_cn428 and end_cn429 and end_cn430 and end_cn431 and end_cn432 and end_cn433 and end_cn434 and end_cn435 and end_cn436 and end_cn437 and end_cn438 and end_cn439 and end_cn440 and end_cn441 and end_cn442 and end_cn443 and end_cn444 and end_cn445 and end_cn446 and end_cn447 and end_cn448 and end_cn449 and end_cn450 and end_cn451 and end_cn452 and end_cn453 and end_cn454 and end_cn455 and end_cn456 and end_cn457 and end_cn458 and end_cn459 and end_cn460 and end_cn461 and end_cn462 and end_cn463 and end_cn464 and end_cn465 and end_cn466 and end_cn467 and end_cn468 and end_cn469 and end_cn470 and end_cn471 and end_cn472 and end_cn473 and end_cn474 and end_cn475 and end_cn476 and end_cn477 and end_cn478 and end_cn479 and end_cn480 and end_cn481 and end_cn482 and end_cn483 and end_cn484 and end_cn485 and end_cn486 and end_cn487 and end_cn488 and end_cn489 and end_cn490 and end_cn491 and end_cn492 and end_cn493 and end_cn494 and end_cn495 and end_cn496 and end_cn497 and end_cn498 and end_cn499 and end_cn500 and end_cn501 and end_cn502 and end_cn503 and end_cn504 and end_cn505 and end_cn506 and end_cn507 and end_cn508 and end_cn509 and end_cn510 and end_cn511 and end_cn512 and end_cn513 and end_cn514 and end_cn515 and end_cn516 and end_cn517 and end_cn518 and end_cn519 and end_cn520 and end_cn521 and end_cn522 and end_cn523 and end_cn524 and end_cn525 and end_cn526 and end_cn527 and end_cn528 and end_cn529 and end_cn530 and end_cn531 and end_cn532 and end_cn533 and end_cn534 and end_cn535 and end_cn536 and end_cn537 and end_cn538 and end_cn539 and end_cn540 and end_cn541 and end_cn542 and end_cn543 and end_cn544 and end_cn545 and end_cn546 and end_cn547 and end_cn548 and end_cn549 and end_cn550 and end_cn551 and end_cn552 and end_cn553 and end_cn554 and end_cn555 and end_cn556 and end_cn557 and end_cn558 and end_cn559 and end_cn560 and end_cn561 and end_cn562 and end_cn563 and end_cn564 and end_cn565 and end_cn566 and end_cn567 and end_cn568 and end_cn569 and end_cn570 and end_cn571 and end_cn572 and end_cn573 and end_cn574 and end_cn575 and end_cn576 and end_cn577 and end_cn578 and end_cn579 and end_cn580 and end_cn581 and end_cn582 and end_cn583 and end_cn584 and end_cn585 and end_cn586 and end_cn587 and end_cn588 and end_cn589 and end_cn590 and end_cn591 and end_cn592 and end_cn593 and end_cn594 and end_cn595 and end_cn596 and end_cn597 and end_cn598 and end_cn599 and end_cn600 and end_cn601 and end_cn602 and end_cn603 and end_cn604 and end_cn605 and end_cn606 and end_cn607 and end_cn608 and end_cn609 and end_cn610 and end_cn611 and end_cn612 and end_cn613 and end_cn614 and end_cn615 and end_cn616 and end_cn617 and end_cn618 and end_cn619 and end_cn620 and end_cn621 and end_cn622 and end_cn623 and end_cn624 and end_cn625 and end_cn626 and end_cn627 and end_cn628 and end_cn629 and end_cn630 and end_cn631 and end_cn632 and end_cn633 and end_cn634 and end_cn635 and end_cn636 and end_cn637 and end_cn638 and end_cn639 and end_cn640 and end_cn641 and end_cn642 and end_cn643 and end_cn644 and end_cn645 and end_cn646 and end_cn647 and end_cn648 and end_cn649 and end_cn650 and end_cn651 and end_cn652 and end_cn653 and end_cn654 and end_cn655 and end_cn656 and end_cn657 and end_cn658 and end_cn659 and end_cn660 and end_cn661 and end_cn662 and end_cn663 and end_cn664 and end_cn665 and end_cn666 and end_cn667 and end_cn668 and end_cn669 and end_cn670 and end_cn671 and end_cn672 and end_cn673 and end_cn674 and end_cn675 and end_cn676 and end_cn677 and end_cn678 and end_cn679 and end_cn680 and end_cn681 and end_cn682 and end_cn683 and end_cn684 and end_cn685 and end_cn686 and end_cn687 and end_cn688 and end_cn689 and end_cn690 and end_cn691 and end_cn692 and end_cn693 and end_cn694 and end_cn695 and end_cn696 and end_cn697 and end_cn698 and end_cn699 and end_cn700 and end_cn701 and end_cn702 and end_cn703 and end_cn704 and end_cn705 and end_cn706 and end_cn707 and end_cn708 and end_cn709 and end_cn710 and end_cn711 and end_cn712 and end_cn713 and end_cn714 and end_cn715 and end_cn716 and end_cn717 and end_cn718 and end_cn719 and end_cn720 and end_cn721 and end_cn722 and end_cn723 and end_cn724 and end_cn725 and end_cn726 and end_cn727 and end_cn728 and end_cn729 and end_cn730 and end_cn731 and end_cn732 and end_cn733 and end_cn734 and end_cn735 and end_cn736 and end_cn737 and end_cn738 and end_cn739 and end_cn740 and end_cn741 and end_cn742 and end_cn743 and end_cn744 and end_cn745 and end_cn746 and end_cn747 and end_cn748 and end_cn749 and end_cn750 and end_cn751 and end_cn752 and end_cn753 and end_cn754 and end_cn755 and end_cn756 and end_cn757 and end_cn758 and end_cn759 and end_cn760 and end_cn761 and end_cn762 and end_cn763 and end_cn764 and end_cn765 and end_cn766 and end_cn767 and end_cn768 and end_cn769 and end_cn770 and end_cn771 and end_cn772 and end_cn773 and end_cn774 and end_cn775 and end_cn776 and end_cn777 and end_cn778 and end_cn779 and end_cn780 and end_cn781 and end_cn782 and end_cn783 and end_cn784 and end_cn785 and end_cn786 and end_cn787 and end_cn788 and end_cn789 and end_cn790 and end_cn791 and end_cn792 and end_cn793 and end_cn794 and end_cn795 and end_cn796 and end_cn797 and end_cn798 and end_cn799 and end_cn800 and end_cn801 and end_cn802 and end_cn803 and end_cn804 and end_cn805 and end_cn806 and end_cn807 and end_cn808 and end_cn809 and end_cn810 and end_cn811 and end_cn812 and end_cn813 and end_cn814 and end_cn815 and end_cn816 and end_cn817 and end_cn818 and end_cn819 and end_cn820 and end_cn821 and end_cn822 and end_cn823 and end_cn824 and end_cn825 and end_cn826 and end_cn827 and end_cn828 and end_cn829 and end_cn830 and end_cn831 and end_cn832 and end_cn833 and end_cn834 and end_cn835 and end_cn836 and end_cn837 and end_cn838 and end_cn839 and end_cn840 and end_cn841 and end_cn842 and end_cn843 and end_cn844 and end_cn845 and end_cn846 and end_cn847 and end_cn848 and end_cn849 and end_cn850 and end_cn851 and end_cn852 and end_cn853 and end_cn854 and end_cn855 and end_cn856 and end_cn857 and end_cn858 and end_cn859 and end_cn860 and end_cn861 and end_cn862 and end_cn863 and end_cn864 and end_cn865 and end_cn866 and end_cn867 and end_cn868 and end_cn869 and end_cn870 and end_cn871 and end_cn872 and end_cn873 and end_cn874 and end_cn875 and end_cn876 and end_cn877 and end_cn878 and end_cn879 and end_cn880 and end_cn881 and end_cn882 and end_cn883 and end_cn884 and end_cn885 and end_cn886 and end_cn887 and end_cn888 and end_cn889 and end_cn890 and end_cn891 and end_cn892 and end_cn893 and end_cn894 and end_cn895 and end_cn896 and end_cn897 and end_cn898 and end_cn899 and end_cn900 and end_cn901 and end_cn902 and end_cn903 and end_cn904 and end_cn905 and end_cn906 and end_cn907 and end_cn908 and end_cn909 and end_cn910 and end_cn911 and end_cn912 and end_cn913 and end_cn914 and end_cn915 and end_cn916 and end_cn917 and end_cn918 and end_cn919 and end_cn920 and end_cn921 and end_cn922 and end_cn923 and end_cn924 and end_cn925 and end_cn926 and end_cn927 and end_cn928 and end_cn929 and end_cn930 and end_cn931 and end_cn932 and end_cn933 and end_cn934 and end_cn935 and end_cn936 and end_cn937 and end_cn938 and end_cn939 and end_cn940 and end_cn941 and end_cn942 and end_cn943 and end_cn944 and end_cn945 and end_cn946 and end_cn947 and end_cn948 and end_cn949 and end_cn950 and end_cn951 and end_cn952 and end_cn953 and end_cn954 and end_cn955 and end_cn956 and end_cn957 and end_cn958 and end_cn959 and end_cn960 and end_cn961 and end_cn962 and end_cn963 and end_cn964 and end_cn965 and end_cn966 and end_cn967 and end_cn968 and end_cn969 and end_cn970 and end_cn971 and end_cn972 and end_cn973 and end_cn974 and end_cn975 and end_cn976 and end_cn977 and end_cn978 and end_cn979 and end_cn980 and end_cn981 and end_cn982 and end_cn983 and end_cn984 and end_cn985 and end_cn986 and end_cn987 and end_cn988 and end_cn989 and end_cn990 and end_cn991 and end_cn992 and end_cn993 and end_cn994 and end_cn995 and end_cn996 and end_cn997 and end_cn998 and end_cn999 and end_cn1000 and end_cn1001 and end_cn1002 and end_cn1003 and end_cn1004 and end_cn1005 and end_cn1006 and end_cn1007 and end_cn1008 and end_cn1009 and end_cn1010 and end_cn1011 and end_cn1012 and end_cn1013 and end_cn1014 and end_cn1015 and end_cn1016 and end_cn1017 and end_cn1018 and end_cn1019 and end_cn1020 and end_cn1021 and end_cn1022 and end_cn1023 and end_cn1024 and end_cn1025 and end_cn1026 and end_cn1027 and end_cn1028 and end_cn1029 and end_cn1030 and end_cn1031 and end_cn1032 and end_cn1033 and end_cn1034 and end_cn1035 and end_cn1036 and end_cn1037 and end_cn1038 and end_cn1039 and end_cn1040 and end_cn1041 and end_cn1042 and end_cn1043 and end_cn1044 and end_cn1045 and end_cn1046 and end_cn1047 and end_cn1048 and end_cn1049 and end_cn1050 and end_cn1051 and end_cn1052 and end_cn1053 and end_cn1054 and end_cn1055 and end_cn1056 and end_cn1057 and end_cn1058 and end_cn1059 and end_cn1060 and end_cn1061 and end_cn1062 and end_cn1063 and end_cn1064 and end_cn1065 and end_cn1066 and end_cn1067 and end_cn1068 and end_cn1069 and end_cn1070 and end_cn1071 and end_cn1072 and end_cn1073 and end_cn1074 and end_cn1075 and end_cn1076 and end_cn1077 and end_cn1078 and end_cn1079 and end_cn1080 and end_cn1081 and end_cn1082 and end_cn1083 and end_cn1084 and end_cn1085 and end_cn1086 and end_cn1087 and end_cn1088 and end_cn1089 and end_cn1090 and end_cn1091 and end_cn1092 and end_cn1093 and end_cn1094 and end_cn1095 and end_cn1096 and end_cn1097 and end_cn1098 and end_cn1099 and end_cn1100 and end_cn1101 and end_cn1102 and end_cn1103 and end_cn1104 and end_cn1105 and end_cn1106 and end_cn1107 and end_cn1108 and end_cn1109 and end_cn1110 and end_cn1111 and end_cn1112 and end_cn1113 and end_cn1114 and end_cn1115 and end_cn1116 and end_cn1117 and end_cn1118 and end_cn1119 and end_cn1120 and end_cn1121 and end_cn1122 and end_cn1123 and end_cn1124 and end_cn1125 and end_cn1126 and end_cn1127 and end_cn1128 and end_cn1129 and end_cn1130 and end_cn1131 and end_cn1132 and end_cn1133 and end_cn1134 and end_cn1135 and end_cn1136 and end_cn1137 and end_cn1138 and end_cn1139 and end_cn1140 and end_cn1141 and end_cn1142 and end_cn1143 and end_cn1144 and end_cn1145 and end_cn1146 and end_cn1147 and end_cn1148 and end_cn1149 and end_cn1150 and end_cn1151 and end_cn1152;
end_vnt<=end_vn1 and end_vn2 and end_vn3 and end_vn4 and end_vn5 and end_vn6 and end_vn7 and end_vn8 and end_vn9 and end_vn10 and end_vn11 and end_vn12 and end_vn13 and end_vn14 and end_vn15 and end_vn16 and end_vn17 and end_vn18 and end_vn19 and end_vn20 and end_vn21 and end_vn22 and end_vn23 and end_vn24 and end_vn25 and end_vn26 and end_vn27 and end_vn28 and end_vn29 and end_vn30 and end_vn31 and end_vn32 and end_vn33 and end_vn34 and end_vn35 and end_vn36 and end_vn37 and end_vn38 and end_vn39 and end_vn40 and end_vn41 and end_vn42 and end_vn43 and end_vn44 and end_vn45 and end_vn46 and end_vn47 and end_vn48 and end_vn49 and end_vn50 and end_vn51 and end_vn52 and end_vn53 and end_vn54 and end_vn55 and end_vn56 and end_vn57 and end_vn58 and end_vn59 and end_vn60 and end_vn61 and end_vn62 and end_vn63 and end_vn64 and end_vn65 and end_vn66 and end_vn67 and end_vn68 and end_vn69 and end_vn70 and end_vn71 and end_vn72 and end_vn73 and end_vn74 and end_vn75 and end_vn76 and end_vn77 and end_vn78 and end_vn79 and end_vn80 and end_vn81 and end_vn82 and end_vn83 and end_vn84 and end_vn85 and end_vn86 and end_vn87 and end_vn88 and end_vn89 and end_vn90 and end_vn91 and end_vn92 and end_vn93 and end_vn94 and end_vn95 and end_vn96 and end_vn97 and end_vn98 and end_vn99 and end_vn100 and end_vn101 and end_vn102 and end_vn103 and end_vn104 and end_vn105 and end_vn106 and end_vn107 and end_vn108 and end_vn109 and end_vn110 and end_vn111 and end_vn112 and end_vn113 and end_vn114 and end_vn115 and end_vn116 and end_vn117 and end_vn118 and end_vn119 and end_vn120 and end_vn121 and end_vn122 and end_vn123 and end_vn124 and end_vn125 and end_vn126 and end_vn127 and end_vn128 and end_vn129 and end_vn130 and end_vn131 and end_vn132 and end_vn133 and end_vn134 and end_vn135 and end_vn136 and end_vn137 and end_vn138 and end_vn139 and end_vn140 and end_vn141 and end_vn142 and end_vn143 and end_vn144 and end_vn145 and end_vn146 and end_vn147 and end_vn148 and end_vn149 and end_vn150 and end_vn151 and end_vn152 and end_vn153 and end_vn154 and end_vn155 and end_vn156 and end_vn157 and end_vn158 and end_vn159 and end_vn160 and end_vn161 and end_vn162 and end_vn163 and end_vn164 and end_vn165 and end_vn166 and end_vn167 and end_vn168 and end_vn169 and end_vn170 and end_vn171 and end_vn172 and end_vn173 and end_vn174 and end_vn175 and end_vn176 and end_vn177 and end_vn178 and end_vn179 and end_vn180 and end_vn181 and end_vn182 and end_vn183 and end_vn184 and end_vn185 and end_vn186 and end_vn187 and end_vn188 and end_vn189 and end_vn190 and end_vn191 and end_vn192 and end_vn193 and end_vn194 and end_vn195 and end_vn196 and end_vn197 and end_vn198 and end_vn199 and end_vn200 and end_vn201 and end_vn202 and end_vn203 and end_vn204 and end_vn205 and end_vn206 and end_vn207 and end_vn208 and end_vn209 and end_vn210 and end_vn211 and end_vn212 and end_vn213 and end_vn214 and end_vn215 and end_vn216 and end_vn217 and end_vn218 and end_vn219 and end_vn220 and end_vn221 and end_vn222 and end_vn223 and end_vn224 and end_vn225 and end_vn226 and end_vn227 and end_vn228 and end_vn229 and end_vn230 and end_vn231 and end_vn232 and end_vn233 and end_vn234 and end_vn235 and end_vn236 and end_vn237 and end_vn238 and end_vn239 and end_vn240 and end_vn241 and end_vn242 and end_vn243 and end_vn244 and end_vn245 and end_vn246 and end_vn247 and end_vn248 and end_vn249 and end_vn250 and end_vn251 and end_vn252 and end_vn253 and end_vn254 and end_vn255 and end_vn256 and end_vn257 and end_vn258 and end_vn259 and end_vn260 and end_vn261 and end_vn262 and end_vn263 and end_vn264 and end_vn265 and end_vn266 and end_vn267 and end_vn268 and end_vn269 and end_vn270 and end_vn271 and end_vn272 and end_vn273 and end_vn274 and end_vn275 and end_vn276 and end_vn277 and end_vn278 and end_vn279 and end_vn280 and end_vn281 and end_vn282 and end_vn283 and end_vn284 and end_vn285 and end_vn286 and end_vn287 and end_vn288 and end_vn289 and end_vn290 and end_vn291 and end_vn292 and end_vn293 and end_vn294 and end_vn295 and end_vn296 and end_vn297 and end_vn298 and end_vn299 and end_vn300 and end_vn301 and end_vn302 and end_vn303 and end_vn304 and end_vn305 and end_vn306 and end_vn307 and end_vn308 and end_vn309 and end_vn310 and end_vn311 and end_vn312 and end_vn313 and end_vn314 and end_vn315 and end_vn316 and end_vn317 and end_vn318 and end_vn319 and end_vn320 and end_vn321 and end_vn322 and end_vn323 and end_vn324 and end_vn325 and end_vn326 and end_vn327 and end_vn328 and end_vn329 and end_vn330 and end_vn331 and end_vn332 and end_vn333 and end_vn334 and end_vn335 and end_vn336 and end_vn337 and end_vn338 and end_vn339 and end_vn340 and end_vn341 and end_vn342 and end_vn343 and end_vn344 and end_vn345 and end_vn346 and end_vn347 and end_vn348 and end_vn349 and end_vn350 and end_vn351 and end_vn352 and end_vn353 and end_vn354 and end_vn355 and end_vn356 and end_vn357 and end_vn358 and end_vn359 and end_vn360 and end_vn361 and end_vn362 and end_vn363 and end_vn364 and end_vn365 and end_vn366 and end_vn367 and end_vn368 and end_vn369 and end_vn370 and end_vn371 and end_vn372 and end_vn373 and end_vn374 and end_vn375 and end_vn376 and end_vn377 and end_vn378 and end_vn379 and end_vn380 and end_vn381 and end_vn382 and end_vn383 and end_vn384 and end_vn385 and end_vn386 and end_vn387 and end_vn388 and end_vn389 and end_vn390 and end_vn391 and end_vn392 and end_vn393 and end_vn394 and end_vn395 and end_vn396 and end_vn397 and end_vn398 and end_vn399 and end_vn400 and end_vn401 and end_vn402 and end_vn403 and end_vn404 and end_vn405 and end_vn406 and end_vn407 and end_vn408 and end_vn409 and end_vn410 and end_vn411 and end_vn412 and end_vn413 and end_vn414 and end_vn415 and end_vn416 and end_vn417 and end_vn418 and end_vn419 and end_vn420 and end_vn421 and end_vn422 and end_vn423 and end_vn424 and end_vn425 and end_vn426 and end_vn427 and end_vn428 and end_vn429 and end_vn430 and end_vn431 and end_vn432 and end_vn433 and end_vn434 and end_vn435 and end_vn436 and end_vn437 and end_vn438 and end_vn439 and end_vn440 and end_vn441 and end_vn442 and end_vn443 and end_vn444 and end_vn445 and end_vn446 and end_vn447 and end_vn448 and end_vn449 and end_vn450 and end_vn451 and end_vn452 and end_vn453 and end_vn454 and end_vn455 and end_vn456 and end_vn457 and end_vn458 and end_vn459 and end_vn460 and end_vn461 and end_vn462 and end_vn463 and end_vn464 and end_vn465 and end_vn466 and end_vn467 and end_vn468 and end_vn469 and end_vn470 and end_vn471 and end_vn472 and end_vn473 and end_vn474 and end_vn475 and end_vn476 and end_vn477 and end_vn478 and end_vn479 and end_vn480 and end_vn481 and end_vn482 and end_vn483 and end_vn484 and end_vn485 and end_vn486 and end_vn487 and end_vn488 and end_vn489 and end_vn490 and end_vn491 and end_vn492 and end_vn493 and end_vn494 and end_vn495 and end_vn496 and end_vn497 and end_vn498 and end_vn499 and end_vn500 and end_vn501 and end_vn502 and end_vn503 and end_vn504 and end_vn505 and end_vn506 and end_vn507 and end_vn508 and end_vn509 and end_vn510 and end_vn511 and end_vn512 and end_vn513 and end_vn514 and end_vn515 and end_vn516 and end_vn517 and end_vn518 and end_vn519 and end_vn520 and end_vn521 and end_vn522 and end_vn523 and end_vn524 and end_vn525 and end_vn526 and end_vn527 and end_vn528 and end_vn529 and end_vn530 and end_vn531 and end_vn532 and end_vn533 and end_vn534 and end_vn535 and end_vn536 and end_vn537 and end_vn538 and end_vn539 and end_vn540 and end_vn541 and end_vn542 and end_vn543 and end_vn544 and end_vn545 and end_vn546 and end_vn547 and end_vn548 and end_vn549 and end_vn550 and end_vn551 and end_vn552 and end_vn553 and end_vn554 and end_vn555 and end_vn556 and end_vn557 and end_vn558 and end_vn559 and end_vn560 and end_vn561 and end_vn562 and end_vn563 and end_vn564 and end_vn565 and end_vn566 and end_vn567 and end_vn568 and end_vn569 and end_vn570 and end_vn571 and end_vn572 and end_vn573 and end_vn574 and end_vn575 and end_vn576 and end_vn577 and end_vn578 and end_vn579 and end_vn580 and end_vn581 and end_vn582 and end_vn583 and end_vn584 and end_vn585 and end_vn586 and end_vn587 and end_vn588 and end_vn589 and end_vn590 and end_vn591 and end_vn592 and end_vn593 and end_vn594 and end_vn595 and end_vn596 and end_vn597 and end_vn598 and end_vn599 and end_vn600 and end_vn601 and end_vn602 and end_vn603 and end_vn604 and end_vn605 and end_vn606 and end_vn607 and end_vn608 and end_vn609 and end_vn610 and end_vn611 and end_vn612 and end_vn613 and end_vn614 and end_vn615 and end_vn616 and end_vn617 and end_vn618 and end_vn619 and end_vn620 and end_vn621 and end_vn622 and end_vn623 and end_vn624 and end_vn625 and end_vn626 and end_vn627 and end_vn628 and end_vn629 and end_vn630 and end_vn631 and end_vn632 and end_vn633 and end_vn634 and end_vn635 and end_vn636 and end_vn637 and end_vn638 and end_vn639 and end_vn640 and end_vn641 and end_vn642 and end_vn643 and end_vn644 and end_vn645 and end_vn646 and end_vn647 and end_vn648 and end_vn649 and end_vn650 and end_vn651 and end_vn652 and end_vn653 and end_vn654 and end_vn655 and end_vn656 and end_vn657 and end_vn658 and end_vn659 and end_vn660 and end_vn661 and end_vn662 and end_vn663 and end_vn664 and end_vn665 and end_vn666 and end_vn667 and end_vn668 and end_vn669 and end_vn670 and end_vn671 and end_vn672 and end_vn673 and end_vn674 and end_vn675 and end_vn676 and end_vn677 and end_vn678 and end_vn679 and end_vn680 and end_vn681 and end_vn682 and end_vn683 and end_vn684 and end_vn685 and end_vn686 and end_vn687 and end_vn688 and end_vn689 and end_vn690 and end_vn691 and end_vn692 and end_vn693 and end_vn694 and end_vn695 and end_vn696 and end_vn697 and end_vn698 and end_vn699 and end_vn700 and end_vn701 and end_vn702 and end_vn703 and end_vn704 and end_vn705 and end_vn706 and end_vn707 and end_vn708 and end_vn709 and end_vn710 and end_vn711 and end_vn712 and end_vn713 and end_vn714 and end_vn715 and end_vn716 and end_vn717 and end_vn718 and end_vn719 and end_vn720 and end_vn721 and end_vn722 and end_vn723 and end_vn724 and end_vn725 and end_vn726 and end_vn727 and end_vn728 and end_vn729 and end_vn730 and end_vn731 and end_vn732 and end_vn733 and end_vn734 and end_vn735 and end_vn736 and end_vn737 and end_vn738 and end_vn739 and end_vn740 and end_vn741 and end_vn742 and end_vn743 and end_vn744 and end_vn745 and end_vn746 and end_vn747 and end_vn748 and end_vn749 and end_vn750 and end_vn751 and end_vn752 and end_vn753 and end_vn754 and end_vn755 and end_vn756 and end_vn757 and end_vn758 and end_vn759 and end_vn760 and end_vn761 and end_vn762 and end_vn763 and end_vn764 and end_vn765 and end_vn766 and end_vn767 and end_vn768 and end_vn769 and end_vn770 and end_vn771 and end_vn772 and end_vn773 and end_vn774 and end_vn775 and end_vn776 and end_vn777 and end_vn778 and end_vn779 and end_vn780 and end_vn781 and end_vn782 and end_vn783 and end_vn784 and end_vn785 and end_vn786 and end_vn787 and end_vn788 and end_vn789 and end_vn790 and end_vn791 and end_vn792 and end_vn793 and end_vn794 and end_vn795 and end_vn796 and end_vn797 and end_vn798 and end_vn799 and end_vn800 and end_vn801 and end_vn802 and end_vn803 and end_vn804 and end_vn805 and end_vn806 and end_vn807 and end_vn808 and end_vn809 and end_vn810 and end_vn811 and end_vn812 and end_vn813 and end_vn814 and end_vn815 and end_vn816 and end_vn817 and end_vn818 and end_vn819 and end_vn820 and end_vn821 and end_vn822 and end_vn823 and end_vn824 and end_vn825 and end_vn826 and end_vn827 and end_vn828 and end_vn829 and end_vn830 and end_vn831 and end_vn832 and end_vn833 and end_vn834 and end_vn835 and end_vn836 and end_vn837 and end_vn838 and end_vn839 and end_vn840 and end_vn841 and end_vn842 and end_vn843 and end_vn844 and end_vn845 and end_vn846 and end_vn847 and end_vn848 and end_vn849 and end_vn850 and end_vn851 and end_vn852 and end_vn853 and end_vn854 and end_vn855 and end_vn856 and end_vn857 and end_vn858 and end_vn859 and end_vn860 and end_vn861 and end_vn862 and end_vn863 and end_vn864 and end_vn865 and end_vn866 and end_vn867 and end_vn868 and end_vn869 and end_vn870 and end_vn871 and end_vn872 and end_vn873 and end_vn874 and end_vn875 and end_vn876 and end_vn877 and end_vn878 and end_vn879 and end_vn880 and end_vn881 and end_vn882 and end_vn883 and end_vn884 and end_vn885 and end_vn886 and end_vn887 and end_vn888 and end_vn889 and end_vn890 and end_vn891 and end_vn892 and end_vn893 and end_vn894 and end_vn895 and end_vn896 and end_vn897 and end_vn898 and end_vn899 and end_vn900 and end_vn901 and end_vn902 and end_vn903 and end_vn904 and end_vn905 and end_vn906 and end_vn907 and end_vn908 and end_vn909 and end_vn910 and end_vn911 and end_vn912 and end_vn913 and end_vn914 and end_vn915 and end_vn916 and end_vn917 and end_vn918 and end_vn919 and end_vn920 and end_vn921 and end_vn922 and end_vn923 and end_vn924 and end_vn925 and end_vn926 and end_vn927 and end_vn928 and end_vn929 and end_vn930 and end_vn931 and end_vn932 and end_vn933 and end_vn934 and end_vn935 and end_vn936 and end_vn937 and end_vn938 and end_vn939 and end_vn940 and end_vn941 and end_vn942 and end_vn943 and end_vn944 and end_vn945 and end_vn946 and end_vn947 and end_vn948 and end_vn949 and end_vn950 and end_vn951 and end_vn952 and end_vn953 and end_vn954 and end_vn955 and end_vn956 and end_vn957 and end_vn958 and end_vn959 and end_vn960 and end_vn961 and end_vn962 and end_vn963 and end_vn964 and end_vn965 and end_vn966 and end_vn967 and end_vn968 and end_vn969 and end_vn970 and end_vn971 and end_vn972 and end_vn973 and end_vn974 and end_vn975 and end_vn976 and end_vn977 and end_vn978 and end_vn979 and end_vn980 and end_vn981 and end_vn982 and end_vn983 and end_vn984 and end_vn985 and end_vn986 and end_vn987 and end_vn988 and end_vn989 and end_vn990 and end_vn991 and end_vn992 and end_vn993 and end_vn994 and end_vn995 and end_vn996 and end_vn997 and end_vn998 and end_vn999 and end_vn1000 and end_vn1001 and end_vn1002 and end_vn1003 and end_vn1004 and end_vn1005 and end_vn1006 and end_vn1007 and end_vn1008 and end_vn1009 and end_vn1010 and end_vn1011 and end_vn1012 and end_vn1013 and end_vn1014 and end_vn1015 and end_vn1016 and end_vn1017 and end_vn1018 and end_vn1019 and end_vn1020 and end_vn1021 and end_vn1022 and end_vn1023 and end_vn1024 and end_vn1025 and end_vn1026 and end_vn1027 and end_vn1028 and end_vn1029 and end_vn1030 and end_vn1031 and end_vn1032 and end_vn1033 and end_vn1034 and end_vn1035 and end_vn1036 and end_vn1037 and end_vn1038 and end_vn1039 and end_vn1040 and end_vn1041 and end_vn1042 and end_vn1043 and end_vn1044 and end_vn1045 and end_vn1046 and end_vn1047 and end_vn1048 and end_vn1049 and end_vn1050 and end_vn1051 and end_vn1052 and end_vn1053 and end_vn1054 and end_vn1055 and end_vn1056 and end_vn1057 and end_vn1058 and end_vn1059 and end_vn1060 and end_vn1061 and end_vn1062 and end_vn1063 and end_vn1064 and end_vn1065 and end_vn1066 and end_vn1067 and end_vn1068 and end_vn1069 and end_vn1070 and end_vn1071 and end_vn1072 and end_vn1073 and end_vn1074 and end_vn1075 and end_vn1076 and end_vn1077 and end_vn1078 and end_vn1079 and end_vn1080 and end_vn1081 and end_vn1082 and end_vn1083 and end_vn1084 and end_vn1085 and end_vn1086 and end_vn1087 and end_vn1088 and end_vn1089 and end_vn1090 and end_vn1091 and end_vn1092 and end_vn1093 and end_vn1094 and end_vn1095 and end_vn1096 and end_vn1097 and end_vn1098 and end_vn1099 and end_vn1100 and end_vn1101 and end_vn1102 and end_vn1103 and end_vn1104 and end_vn1105 and end_vn1106 and end_vn1107 and end_vn1108 and end_vn1109 and end_vn1110 and end_vn1111 and end_vn1112 and end_vn1113 and end_vn1114 and end_vn1115 and end_vn1116 and end_vn1117 and end_vn1118 and end_vn1119 and end_vn1120 and end_vn1121 and end_vn1122 and end_vn1123 and end_vn1124 and end_vn1125 and end_vn1126 and end_vn1127 and end_vn1128 and end_vn1129 and end_vn1130 and end_vn1131 and end_vn1132 and end_vn1133 and end_vn1134 and end_vn1135 and end_vn1136 and end_vn1137 and end_vn1138 and end_vn1139 and end_vn1140 and end_vn1141 and end_vn1142 and end_vn1143 and end_vn1144 and end_vn1145 and end_vn1146 and end_vn1147 and end_vn1148 and end_vn1149 and end_vn1150 and end_vn1151 and end_vn1152 and end_vn1153 and end_vn1154 and end_vn1155 and end_vn1156 and end_vn1157 and end_vn1158 and end_vn1159 and end_vn1160 and end_vn1161 and end_vn1162 and end_vn1163 and end_vn1164 and end_vn1165 and end_vn1166 and end_vn1167 and end_vn1168 and end_vn1169 and end_vn1170 and end_vn1171 and end_vn1172 and end_vn1173 and end_vn1174 and end_vn1175 and end_vn1176 and end_vn1177 and end_vn1178 and end_vn1179 and end_vn1180 and end_vn1181 and end_vn1182 and end_vn1183 and end_vn1184 and end_vn1185 and end_vn1186 and end_vn1187 and end_vn1188 and end_vn1189 and end_vn1190 and end_vn1191 and end_vn1192 and end_vn1193 and end_vn1194 and end_vn1195 and end_vn1196 and end_vn1197 and end_vn1198 and end_vn1199 and end_vn1200 and end_vn1201 and end_vn1202 and end_vn1203 and end_vn1204 and end_vn1205 and end_vn1206 and end_vn1207 and end_vn1208 and end_vn1209 and end_vn1210 and end_vn1211 and end_vn1212 and end_vn1213 and end_vn1214 and end_vn1215 and end_vn1216 and end_vn1217 and end_vn1218 and end_vn1219 and end_vn1220 and end_vn1221 and end_vn1222 and end_vn1223 and end_vn1224 and end_vn1225 and end_vn1226 and end_vn1227 and end_vn1228 and end_vn1229 and end_vn1230 and end_vn1231 and end_vn1232 and end_vn1233 and end_vn1234 and end_vn1235 and end_vn1236 and end_vn1237 and end_vn1238 and end_vn1239 and end_vn1240 and end_vn1241 and end_vn1242 and end_vn1243 and end_vn1244 and end_vn1245 and end_vn1246 and end_vn1247 and end_vn1248 and end_vn1249 and end_vn1250 and end_vn1251 and end_vn1252 and end_vn1253 and end_vn1254 and end_vn1255 and end_vn1256 and end_vn1257 and end_vn1258 and end_vn1259 and end_vn1260 and end_vn1261 and end_vn1262 and end_vn1263 and end_vn1264 and end_vn1265 and end_vn1266 and end_vn1267 and end_vn1268 and end_vn1269 and end_vn1270 and end_vn1271 and end_vn1272 and end_vn1273 and end_vn1274 and end_vn1275 and end_vn1276 and end_vn1277 and end_vn1278 and end_vn1279 and end_vn1280 and end_vn1281 and end_vn1282 and end_vn1283 and end_vn1284 and end_vn1285 and end_vn1286 and end_vn1287 and end_vn1288 and end_vn1289 and end_vn1290 and end_vn1291 and end_vn1292 and end_vn1293 and end_vn1294 and end_vn1295 and end_vn1296 and end_vn1297 and end_vn1298 and end_vn1299 and end_vn1300 and end_vn1301 and end_vn1302 and end_vn1303 and end_vn1304 and end_vn1305 and end_vn1306 and end_vn1307 and end_vn1308 and end_vn1309 and end_vn1310 and end_vn1311 and end_vn1312 and end_vn1313 and end_vn1314 and end_vn1315 and end_vn1316 and end_vn1317 and end_vn1318 and end_vn1319 and end_vn1320 and end_vn1321 and end_vn1322 and end_vn1323 and end_vn1324 and end_vn1325 and end_vn1326 and end_vn1327 and end_vn1328 and end_vn1329 and end_vn1330 and end_vn1331 and end_vn1332 and end_vn1333 and end_vn1334 and end_vn1335 and end_vn1336 and end_vn1337 and end_vn1338 and end_vn1339 and end_vn1340 and end_vn1341 and end_vn1342 and end_vn1343 and end_vn1344 and end_vn1345 and end_vn1346 and end_vn1347 and end_vn1348 and end_vn1349 and end_vn1350 and end_vn1351 and end_vn1352 and end_vn1353 and end_vn1354 and end_vn1355 and end_vn1356 and end_vn1357 and end_vn1358 and end_vn1359 and end_vn1360 and end_vn1361 and end_vn1362 and end_vn1363 and end_vn1364 and end_vn1365 and end_vn1366 and end_vn1367 and end_vn1368 and end_vn1369 and end_vn1370 and end_vn1371 and end_vn1372 and end_vn1373 and end_vn1374 and end_vn1375 and end_vn1376 and end_vn1377 and end_vn1378 and end_vn1379 and end_vn1380 and end_vn1381 and end_vn1382 and end_vn1383 and end_vn1384 and end_vn1385 and end_vn1386 and end_vn1387 and end_vn1388 and end_vn1389 and end_vn1390 and end_vn1391 and end_vn1392 and end_vn1393 and end_vn1394 and end_vn1395 and end_vn1396 and end_vn1397 and end_vn1398 and end_vn1399 and end_vn1400 and end_vn1401 and end_vn1402 and end_vn1403 and end_vn1404 and end_vn1405 and end_vn1406 and end_vn1407 and end_vn1408 and end_vn1409 and end_vn1410 and end_vn1411 and end_vn1412 and end_vn1413 and end_vn1414 and end_vn1415 and end_vn1416 and end_vn1417 and end_vn1418 and end_vn1419 and end_vn1420 and end_vn1421 and end_vn1422 and end_vn1423 and end_vn1424 and end_vn1425 and end_vn1426 and end_vn1427 and end_vn1428 and end_vn1429 and end_vn1430 and end_vn1431 and end_vn1432 and end_vn1433 and end_vn1434 and end_vn1435 and end_vn1436 and end_vn1437 and end_vn1438 and end_vn1439 and end_vn1440 and end_vn1441 and end_vn1442 and end_vn1443 and end_vn1444 and end_vn1445 and end_vn1446 and end_vn1447 and end_vn1448 and end_vn1449 and end_vn1450 and end_vn1451 and end_vn1452 and end_vn1453 and end_vn1454 and end_vn1455 and end_vn1456 and end_vn1457 and end_vn1458 and end_vn1459 and end_vn1460 and end_vn1461 and end_vn1462 and end_vn1463 and end_vn1464 and end_vn1465 and end_vn1466 and end_vn1467 and end_vn1468 and end_vn1469 and end_vn1470 and end_vn1471 and end_vn1472 and end_vn1473 and end_vn1474 and end_vn1475 and end_vn1476 and end_vn1477 and end_vn1478 and end_vn1479 and end_vn1480 and end_vn1481 and end_vn1482 and end_vn1483 and end_vn1484 and end_vn1485 and end_vn1486 and end_vn1487 and end_vn1488 and end_vn1489 and end_vn1490 and end_vn1491 and end_vn1492 and end_vn1493 and end_vn1494 and end_vn1495 and end_vn1496 and end_vn1497 and end_vn1498 and end_vn1499 and end_vn1500 and end_vn1501 and end_vn1502 and end_vn1503 and end_vn1504 and end_vn1505 and end_vn1506 and end_vn1507 and end_vn1508 and end_vn1509 and end_vn1510 and end_vn1511 and end_vn1512 and end_vn1513 and end_vn1514 and end_vn1515 and end_vn1516 and end_vn1517 and end_vn1518 and end_vn1519 and end_vn1520 and end_vn1521 and end_vn1522 and end_vn1523 and end_vn1524 and end_vn1525 and end_vn1526 and end_vn1527 and end_vn1528 and end_vn1529 and end_vn1530 and end_vn1531 and end_vn1532 and end_vn1533 and end_vn1534 and end_vn1535 and end_vn1536 and end_vn1537 and end_vn1538 and end_vn1539 and end_vn1540 and end_vn1541 and end_vn1542 and end_vn1543 and end_vn1544 and end_vn1545 and end_vn1546 and end_vn1547 and end_vn1548 and end_vn1549 and end_vn1550 and end_vn1551 and end_vn1552 and end_vn1553 and end_vn1554 and end_vn1555 and end_vn1556 and end_vn1557 and end_vn1558 and end_vn1559 and end_vn1560 and end_vn1561 and end_vn1562 and end_vn1563 and end_vn1564 and end_vn1565 and end_vn1566 and end_vn1567 and end_vn1568 and end_vn1569 and end_vn1570 and end_vn1571 and end_vn1572 and end_vn1573 and end_vn1574 and end_vn1575 and end_vn1576 and end_vn1577 and end_vn1578 and end_vn1579 and end_vn1580 and end_vn1581 and end_vn1582 and end_vn1583 and end_vn1584 and end_vn1585 and end_vn1586 and end_vn1587 and end_vn1588 and end_vn1589 and end_vn1590 and end_vn1591 and end_vn1592 and end_vn1593 and end_vn1594 and end_vn1595 and end_vn1596 and end_vn1597 and end_vn1598 and end_vn1599 and end_vn1600 and end_vn1601 and end_vn1602 and end_vn1603 and end_vn1604 and end_vn1605 and end_vn1606 and end_vn1607 and end_vn1608 and end_vn1609 and end_vn1610 and end_vn1611 and end_vn1612 and end_vn1613 and end_vn1614 and end_vn1615 and end_vn1616 and end_vn1617 and end_vn1618 and end_vn1619 and end_vn1620 and end_vn1621 and end_vn1622 and end_vn1623 and end_vn1624 and end_vn1625 and end_vn1626 and end_vn1627 and end_vn1628 and end_vn1629 and end_vn1630 and end_vn1631 and end_vn1632 and end_vn1633 and end_vn1634 and end_vn1635 and end_vn1636 and end_vn1637 and end_vn1638 and end_vn1639 and end_vn1640 and end_vn1641 and end_vn1642 and end_vn1643 and end_vn1644 and end_vn1645 and end_vn1646 and end_vn1647 and end_vn1648 and end_vn1649 and end_vn1650 and end_vn1651 and end_vn1652 and end_vn1653 and end_vn1654 and end_vn1655 and end_vn1656 and end_vn1657 and end_vn1658 and end_vn1659 and end_vn1660 and end_vn1661 and end_vn1662 and end_vn1663 and end_vn1664 and end_vn1665 and end_vn1666 and end_vn1667 and end_vn1668 and end_vn1669 and end_vn1670 and end_vn1671 and end_vn1672 and end_vn1673 and end_vn1674 and end_vn1675 and end_vn1676 and end_vn1677 and end_vn1678 and end_vn1679 and end_vn1680 and end_vn1681 and end_vn1682 and end_vn1683 and end_vn1684 and end_vn1685 and end_vn1686 and end_vn1687 and end_vn1688 and end_vn1689 and end_vn1690 and end_vn1691 and end_vn1692 and end_vn1693 and end_vn1694 and end_vn1695 and end_vn1696 and end_vn1697 and end_vn1698 and end_vn1699 and end_vn1700 and end_vn1701 and end_vn1702 and end_vn1703 and end_vn1704 and end_vn1705 and end_vn1706 and end_vn1707 and end_vn1708 and end_vn1709 and end_vn1710 and end_vn1711 and end_vn1712 and end_vn1713 and end_vn1714 and end_vn1715 and end_vn1716 and end_vn1717 and end_vn1718 and end_vn1719 and end_vn1720 and end_vn1721 and end_vn1722 and end_vn1723 and end_vn1724 and end_vn1725 and end_vn1726 and end_vn1727 and end_vn1728 and end_vn1729 and end_vn1730 and end_vn1731 and end_vn1732 and end_vn1733 and end_vn1734 and end_vn1735 and end_vn1736 and end_vn1737 and end_vn1738 and end_vn1739 and end_vn1740 and end_vn1741 and end_vn1742 and end_vn1743 and end_vn1744 and end_vn1745 and end_vn1746 and end_vn1747 and end_vn1748 and end_vn1749 and end_vn1750 and end_vn1751 and end_vn1752 and end_vn1753 and end_vn1754 and end_vn1755 and end_vn1756 and end_vn1757 and end_vn1758 and end_vn1759 and end_vn1760 and end_vn1761 and end_vn1762 and end_vn1763 and end_vn1764 and end_vn1765 and end_vn1766 and end_vn1767 and end_vn1768 and end_vn1769 and end_vn1770 and end_vn1771 and end_vn1772 and end_vn1773 and end_vn1774 and end_vn1775 and end_vn1776 and end_vn1777 and end_vn1778 and end_vn1779 and end_vn1780 and end_vn1781 and end_vn1782 and end_vn1783 and end_vn1784 and end_vn1785 and end_vn1786 and end_vn1787 and end_vn1788 and end_vn1789 and end_vn1790 and end_vn1791 and end_vn1792 and end_vn1793 and end_vn1794 and end_vn1795 and end_vn1796 and end_vn1797 and end_vn1798 and end_vn1799 and end_vn1800 and end_vn1801 and end_vn1802 and end_vn1803 and end_vn1804 and end_vn1805 and end_vn1806 and end_vn1807 and end_vn1808 and end_vn1809 and end_vn1810 and end_vn1811 and end_vn1812 and end_vn1813 and end_vn1814 and end_vn1815 and end_vn1816 and end_vn1817 and end_vn1818 and end_vn1819 and end_vn1820 and end_vn1821 and end_vn1822 and end_vn1823 and end_vn1824 and end_vn1825 and end_vn1826 and end_vn1827 and end_vn1828 and end_vn1829 and end_vn1830 and end_vn1831 and end_vn1832 and end_vn1833 and end_vn1834 and end_vn1835 and end_vn1836 and end_vn1837 and end_vn1838 and end_vn1839 and end_vn1840 and end_vn1841 and end_vn1842 and end_vn1843 and end_vn1844 and end_vn1845 and end_vn1846 and end_vn1847 and end_vn1848 and end_vn1849 and end_vn1850 and end_vn1851 and end_vn1852 and end_vn1853 and end_vn1854 and end_vn1855 and end_vn1856 and end_vn1857 and end_vn1858 and end_vn1859 and end_vn1860 and end_vn1861 and end_vn1862 and end_vn1863 and end_vn1864 and end_vn1865 and end_vn1866 and end_vn1867 and end_vn1868 and end_vn1869 and end_vn1870 and end_vn1871 and end_vn1872 and end_vn1873 and end_vn1874 and end_vn1875 and end_vn1876 and end_vn1877 and end_vn1878 and end_vn1879 and end_vn1880 and end_vn1881 and end_vn1882 and end_vn1883 and end_vn1884 and end_vn1885 and end_vn1886 and end_vn1887 and end_vn1888 and end_vn1889 and end_vn1890 and end_vn1891 and end_vn1892 and end_vn1893 and end_vn1894 and end_vn1895 and end_vn1896 and end_vn1897 and end_vn1898 and end_vn1899 and end_vn1900 and end_vn1901 and end_vn1902 and end_vn1903 and end_vn1904 and end_vn1905 and end_vn1906 and end_vn1907 and end_vn1908 and end_vn1909 and end_vn1910 and end_vn1911 and end_vn1912 and end_vn1913 and end_vn1914 and end_vn1915 and end_vn1916 and end_vn1917 and end_vn1918 and end_vn1919 and end_vn1920 and end_vn1921 and end_vn1922 and end_vn1923 and end_vn1924 and end_vn1925 and end_vn1926 and end_vn1927 and end_vn1928 and end_vn1929 and end_vn1930 and end_vn1931 and end_vn1932 and end_vn1933 and end_vn1934 and end_vn1935 and end_vn1936 and end_vn1937 and end_vn1938 and end_vn1939 and end_vn1940 and end_vn1941 and end_vn1942 and end_vn1943 and end_vn1944 and end_vn1945 and end_vn1946 and end_vn1947 and end_vn1948 and end_vn1949 and end_vn1950 and end_vn1951 and end_vn1952 and end_vn1953 and end_vn1954 and end_vn1955 and end_vn1956 and end_vn1957 and end_vn1958 and end_vn1959 and end_vn1960 and end_vn1961 and end_vn1962 and end_vn1963 and end_vn1964 and end_vn1965 and end_vn1966 and end_vn1967 and end_vn1968 and end_vn1969 and end_vn1970 and end_vn1971 and end_vn1972 and end_vn1973 and end_vn1974 and end_vn1975 and end_vn1976 and end_vn1977 and end_vn1978 and end_vn1979 and end_vn1980 and end_vn1981 and end_vn1982 and end_vn1983 and end_vn1984 and end_vn1985 and end_vn1986 and end_vn1987 and end_vn1988 and end_vn1989 and end_vn1990 and end_vn1991 and end_vn1992 and end_vn1993 and end_vn1994 and end_vn1995 and end_vn1996 and end_vn1997 and end_vn1998 and end_vn1999 and end_vn2000 and end_vn2001 and end_vn2002 and end_vn2003 and end_vn2004 and end_vn2005 and end_vn2006 and end_vn2007 and end_vn2008 and end_vn2009 and end_vn2010 and end_vn2011 and end_vn2012 and end_vn2013 and end_vn2014 and end_vn2015 and end_vn2016 and end_vn2017 and end_vn2018 and end_vn2019 and end_vn2020 and end_vn2021 and end_vn2022 and end_vn2023 and end_vn2024 and end_vn2025 and end_vn2026 and end_vn2027 and end_vn2028 and end_vn2029 and end_vn2030 and end_vn2031 and end_vn2032 and end_vn2033 and end_vn2034 and end_vn2035 and end_vn2036 and end_vn2037 and end_vn2038 and end_vn2039 and end_vn2040 and end_vn2041 and end_vn2042 and end_vn2043 and end_vn2044 and end_vn2045 and end_vn2046 and end_vn2047 and end_vn2048 and end_vn2049 and end_vn2050 and end_vn2051 and end_vn2052 and end_vn2053 and end_vn2054 and end_vn2055 and end_vn2056 and end_vn2057 and end_vn2058 and end_vn2059 and end_vn2060 and end_vn2061 and end_vn2062 and end_vn2063 and end_vn2064 and end_vn2065 and end_vn2066 and end_vn2067 and end_vn2068 and end_vn2069 and end_vn2070 and end_vn2071 and end_vn2072 and end_vn2073 and end_vn2074 and end_vn2075 and end_vn2076 and end_vn2077 and end_vn2078 and end_vn2079 and end_vn2080 and end_vn2081 and end_vn2082 and end_vn2083 and end_vn2084 and end_vn2085 and end_vn2086 and end_vn2087 and end_vn2088 and end_vn2089 and end_vn2090 and end_vn2091 and end_vn2092 and end_vn2093 and end_vn2094 and end_vn2095 and end_vn2096 and end_vn2097 and end_vn2098 and end_vn2099 and end_vn2100 and end_vn2101 and end_vn2102 and end_vn2103 and end_vn2104 and end_vn2105 and end_vn2106 and end_vn2107 and end_vn2108 and end_vn2109 and end_vn2110 and end_vn2111 and end_vn2112 and end_vn2113 and end_vn2114 and end_vn2115 and end_vn2116 and end_vn2117 and end_vn2118 and end_vn2119 and end_vn2120 and end_vn2121 and end_vn2122 and end_vn2123 and end_vn2124 and end_vn2125 and end_vn2126 and end_vn2127 and end_vn2128 and end_vn2129 and end_vn2130 and end_vn2131 and end_vn2132 and end_vn2133 and end_vn2134 and end_vn2135 and end_vn2136 and end_vn2137 and end_vn2138 and end_vn2139 and end_vn2140 and end_vn2141 and end_vn2142 and end_vn2143 and end_vn2144 and end_vn2145 and end_vn2146 and end_vn2147 and end_vn2148 and end_vn2149 and end_vn2150 and end_vn2151 and end_vn2152 and end_vn2153 and end_vn2154 and end_vn2155 and end_vn2156 and end_vn2157 and end_vn2158 and end_vn2159 and end_vn2160 and end_vn2161 and end_vn2162 and end_vn2163 and end_vn2164 and end_vn2165 and end_vn2166 and end_vn2167 and end_vn2168 and end_vn2169 and end_vn2170 and end_vn2171 and end_vn2172 and end_vn2173 and end_vn2174 and end_vn2175 and end_vn2176 and end_vn2177 and end_vn2178 and end_vn2179 and end_vn2180 and end_vn2181 and end_vn2182 and end_vn2183 and end_vn2184 and end_vn2185 and end_vn2186 and end_vn2187 and end_vn2188 and end_vn2189 and end_vn2190 and end_vn2191 and end_vn2192 and end_vn2193 and end_vn2194 and end_vn2195 and end_vn2196 and end_vn2197 and end_vn2198 and end_vn2199 and end_vn2200 and end_vn2201 and end_vn2202 and end_vn2203 and end_vn2204 and end_vn2205 and end_vn2206 and end_vn2207 and end_vn2208 and end_vn2209 and end_vn2210 and end_vn2211 and end_vn2212 and end_vn2213 and end_vn2214 and end_vn2215 and end_vn2216 and end_vn2217 and end_vn2218 and end_vn2219 and end_vn2220 and end_vn2221 and end_vn2222 and end_vn2223 and end_vn2224 and end_vn2225 and end_vn2226 and end_vn2227 and end_vn2228 and end_vn2229 and end_vn2230 and end_vn2231 and end_vn2232 and end_vn2233 and end_vn2234 and end_vn2235 and end_vn2236 and end_vn2237 and end_vn2238 and end_vn2239 and end_vn2240 and end_vn2241 and end_vn2242 and end_vn2243 and end_vn2244 and end_vn2245 and end_vn2246 and end_vn2247 and end_vn2248 and end_vn2249 and end_vn2250 and end_vn2251 and end_vn2252 and end_vn2253 and end_vn2254 and end_vn2255 and end_vn2256 and end_vn2257 and end_vn2258 and end_vn2259 and end_vn2260 and end_vn2261 and end_vn2262 and end_vn2263 and end_vn2264 and end_vn2265 and end_vn2266 and end_vn2267 and end_vn2268 and end_vn2269 and end_vn2270 and end_vn2271 and end_vn2272 and end_vn2273 and end_vn2274 and end_vn2275 and end_vn2276 and end_vn2277 and end_vn2278 and end_vn2279 and end_vn2280 and end_vn2281 and end_vn2282 and end_vn2283 and end_vn2284 and end_vn2285 and end_vn2286 and end_vn2287 and end_vn2288 and end_vn2289 and end_vn2290 and end_vn2291 and end_vn2292 and end_vn2293 and end_vn2294 and end_vn2295 and end_vn2296 and end_vn2297 and end_vn2298 and end_vn2299 and end_vn2300 and end_vn2301 and end_vn2302 and end_vn2303 and end_vn2304;
out1<=SI1;
out2<=SI2;
out3<=SI3;
out4<=SI4;
out5<=SI5;
out6<=SI6;
out7<=SI7;
out8<=SI8;
out9<=SI9;
out10<=SI10;
out11<=SI11;
out12<=SI12;
out13<=SI13;
out14<=SI14;
out15<=SI15;
out16<=SI16;
out17<=SI17;
out18<=SI18;
out19<=SI19;
out20<=SI20;
out21<=SI21;
out22<=SI22;
out23<=SI23;
out24<=SI24;
out25<=SI25;
out26<=SI26;
out27<=SI27;
out28<=SI28;
out29<=SI29;
out30<=SI30;
out31<=SI31;
out32<=SI32;
out33<=SI33;
out34<=SI34;
out35<=SI35;
out36<=SI36;
out37<=SI37;
out38<=SI38;
out39<=SI39;
out40<=SI40;
out41<=SI41;
out42<=SI42;
out43<=SI43;
out44<=SI44;
out45<=SI45;
out46<=SI46;
out47<=SI47;
out48<=SI48;
out49<=SI49;
out50<=SI50;
out51<=SI51;
out52<=SI52;
out53<=SI53;
out54<=SI54;
out55<=SI55;
out56<=SI56;
out57<=SI57;
out58<=SI58;
out59<=SI59;
out60<=SI60;
out61<=SI61;
out62<=SI62;
out63<=SI63;
out64<=SI64;
out65<=SI65;
out66<=SI66;
out67<=SI67;
out68<=SI68;
out69<=SI69;
out70<=SI70;
out71<=SI71;
out72<=SI72;
out73<=SI73;
out74<=SI74;
out75<=SI75;
out76<=SI76;
out77<=SI77;
out78<=SI78;
out79<=SI79;
out80<=SI80;
out81<=SI81;
out82<=SI82;
out83<=SI83;
out84<=SI84;
out85<=SI85;
out86<=SI86;
out87<=SI87;
out88<=SI88;
out89<=SI89;
out90<=SI90;
out91<=SI91;
out92<=SI92;
out93<=SI93;
out94<=SI94;
out95<=SI95;
out96<=SI96;
out97<=SI97;
out98<=SI98;
out99<=SI99;
out100<=SI100;
out101<=SI101;
out102<=SI102;
out103<=SI103;
out104<=SI104;
out105<=SI105;
out106<=SI106;
out107<=SI107;
out108<=SI108;
out109<=SI109;
out110<=SI110;
out111<=SI111;
out112<=SI112;
out113<=SI113;
out114<=SI114;
out115<=SI115;
out116<=SI116;
out117<=SI117;
out118<=SI118;
out119<=SI119;
out120<=SI120;
out121<=SI121;
out122<=SI122;
out123<=SI123;
out124<=SI124;
out125<=SI125;
out126<=SI126;
out127<=SI127;
out128<=SI128;
out129<=SI129;
out130<=SI130;
out131<=SI131;
out132<=SI132;
out133<=SI133;
out134<=SI134;
out135<=SI135;
out136<=SI136;
out137<=SI137;
out138<=SI138;
out139<=SI139;
out140<=SI140;
out141<=SI141;
out142<=SI142;
out143<=SI143;
out144<=SI144;
out145<=SI145;
out146<=SI146;
out147<=SI147;
out148<=SI148;
out149<=SI149;
out150<=SI150;
out151<=SI151;
out152<=SI152;
out153<=SI153;
out154<=SI154;
out155<=SI155;
out156<=SI156;
out157<=SI157;
out158<=SI158;
out159<=SI159;
out160<=SI160;
out161<=SI161;
out162<=SI162;
out163<=SI163;
out164<=SI164;
out165<=SI165;
out166<=SI166;
out167<=SI167;
out168<=SI168;
out169<=SI169;
out170<=SI170;
out171<=SI171;
out172<=SI172;
out173<=SI173;
out174<=SI174;
out175<=SI175;
out176<=SI176;
out177<=SI177;
out178<=SI178;
out179<=SI179;
out180<=SI180;
out181<=SI181;
out182<=SI182;
out183<=SI183;
out184<=SI184;
out185<=SI185;
out186<=SI186;
out187<=SI187;
out188<=SI188;
out189<=SI189;
out190<=SI190;
out191<=SI191;
out192<=SI192;
out193<=SI193;
out194<=SI194;
out195<=SI195;
out196<=SI196;
out197<=SI197;
out198<=SI198;
out199<=SI199;
out200<=SI200;
out201<=SI201;
out202<=SI202;
out203<=SI203;
out204<=SI204;
out205<=SI205;
out206<=SI206;
out207<=SI207;
out208<=SI208;
out209<=SI209;
out210<=SI210;
out211<=SI211;
out212<=SI212;
out213<=SI213;
out214<=SI214;
out215<=SI215;
out216<=SI216;
out217<=SI217;
out218<=SI218;
out219<=SI219;
out220<=SI220;
out221<=SI221;
out222<=SI222;
out223<=SI223;
out224<=SI224;
out225<=SI225;
out226<=SI226;
out227<=SI227;
out228<=SI228;
out229<=SI229;
out230<=SI230;
out231<=SI231;
out232<=SI232;
out233<=SI233;
out234<=SI234;
out235<=SI235;
out236<=SI236;
out237<=SI237;
out238<=SI238;
out239<=SI239;
out240<=SI240;
out241<=SI241;
out242<=SI242;
out243<=SI243;
out244<=SI244;
out245<=SI245;
out246<=SI246;
out247<=SI247;
out248<=SI248;
out249<=SI249;
out250<=SI250;
out251<=SI251;
out252<=SI252;
out253<=SI253;
out254<=SI254;
out255<=SI255;
out256<=SI256;
out257<=SI257;
out258<=SI258;
out259<=SI259;
out260<=SI260;
out261<=SI261;
out262<=SI262;
out263<=SI263;
out264<=SI264;
out265<=SI265;
out266<=SI266;
out267<=SI267;
out268<=SI268;
out269<=SI269;
out270<=SI270;
out271<=SI271;
out272<=SI272;
out273<=SI273;
out274<=SI274;
out275<=SI275;
out276<=SI276;
out277<=SI277;
out278<=SI278;
out279<=SI279;
out280<=SI280;
out281<=SI281;
out282<=SI282;
out283<=SI283;
out284<=SI284;
out285<=SI285;
out286<=SI286;
out287<=SI287;
out288<=SI288;
out289<=SI289;
out290<=SI290;
out291<=SI291;
out292<=SI292;
out293<=SI293;
out294<=SI294;
out295<=SI295;
out296<=SI296;
out297<=SI297;
out298<=SI298;
out299<=SI299;
out300<=SI300;
out301<=SI301;
out302<=SI302;
out303<=SI303;
out304<=SI304;
out305<=SI305;
out306<=SI306;
out307<=SI307;
out308<=SI308;
out309<=SI309;
out310<=SI310;
out311<=SI311;
out312<=SI312;
out313<=SI313;
out314<=SI314;
out315<=SI315;
out316<=SI316;
out317<=SI317;
out318<=SI318;
out319<=SI319;
out320<=SI320;
out321<=SI321;
out322<=SI322;
out323<=SI323;
out324<=SI324;
out325<=SI325;
out326<=SI326;
out327<=SI327;
out328<=SI328;
out329<=SI329;
out330<=SI330;
out331<=SI331;
out332<=SI332;
out333<=SI333;
out334<=SI334;
out335<=SI335;
out336<=SI336;
out337<=SI337;
out338<=SI338;
out339<=SI339;
out340<=SI340;
out341<=SI341;
out342<=SI342;
out343<=SI343;
out344<=SI344;
out345<=SI345;
out346<=SI346;
out347<=SI347;
out348<=SI348;
out349<=SI349;
out350<=SI350;
out351<=SI351;
out352<=SI352;
out353<=SI353;
out354<=SI354;
out355<=SI355;
out356<=SI356;
out357<=SI357;
out358<=SI358;
out359<=SI359;
out360<=SI360;
out361<=SI361;
out362<=SI362;
out363<=SI363;
out364<=SI364;
out365<=SI365;
out366<=SI366;
out367<=SI367;
out368<=SI368;
out369<=SI369;
out370<=SI370;
out371<=SI371;
out372<=SI372;
out373<=SI373;
out374<=SI374;
out375<=SI375;
out376<=SI376;
out377<=SI377;
out378<=SI378;
out379<=SI379;
out380<=SI380;
out381<=SI381;
out382<=SI382;
out383<=SI383;
out384<=SI384;
out385<=SI385;
out386<=SI386;
out387<=SI387;
out388<=SI388;
out389<=SI389;
out390<=SI390;
out391<=SI391;
out392<=SI392;
out393<=SI393;
out394<=SI394;
out395<=SI395;
out396<=SI396;
out397<=SI397;
out398<=SI398;
out399<=SI399;
out400<=SI400;
out401<=SI401;
out402<=SI402;
out403<=SI403;
out404<=SI404;
out405<=SI405;
out406<=SI406;
out407<=SI407;
out408<=SI408;
out409<=SI409;
out410<=SI410;
out411<=SI411;
out412<=SI412;
out413<=SI413;
out414<=SI414;
out415<=SI415;
out416<=SI416;
out417<=SI417;
out418<=SI418;
out419<=SI419;
out420<=SI420;
out421<=SI421;
out422<=SI422;
out423<=SI423;
out424<=SI424;
out425<=SI425;
out426<=SI426;
out427<=SI427;
out428<=SI428;
out429<=SI429;
out430<=SI430;
out431<=SI431;
out432<=SI432;
out433<=SI433;
out434<=SI434;
out435<=SI435;
out436<=SI436;
out437<=SI437;
out438<=SI438;
out439<=SI439;
out440<=SI440;
out441<=SI441;
out442<=SI442;
out443<=SI443;
out444<=SI444;
out445<=SI445;
out446<=SI446;
out447<=SI447;
out448<=SI448;
out449<=SI449;
out450<=SI450;
out451<=SI451;
out452<=SI452;
out453<=SI453;
out454<=SI454;
out455<=SI455;
out456<=SI456;
out457<=SI457;
out458<=SI458;
out459<=SI459;
out460<=SI460;
out461<=SI461;
out462<=SI462;
out463<=SI463;
out464<=SI464;
out465<=SI465;
out466<=SI466;
out467<=SI467;
out468<=SI468;
out469<=SI469;
out470<=SI470;
out471<=SI471;
out472<=SI472;
out473<=SI473;
out474<=SI474;
out475<=SI475;
out476<=SI476;
out477<=SI477;
out478<=SI478;
out479<=SI479;
out480<=SI480;
out481<=SI481;
out482<=SI482;
out483<=SI483;
out484<=SI484;
out485<=SI485;
out486<=SI486;
out487<=SI487;
out488<=SI488;
out489<=SI489;
out490<=SI490;
out491<=SI491;
out492<=SI492;
out493<=SI493;
out494<=SI494;
out495<=SI495;
out496<=SI496;
out497<=SI497;
out498<=SI498;
out499<=SI499;
out500<=SI500;
out501<=SI501;
out502<=SI502;
out503<=SI503;
out504<=SI504;
out505<=SI505;
out506<=SI506;
out507<=SI507;
out508<=SI508;
out509<=SI509;
out510<=SI510;
out511<=SI511;
out512<=SI512;
out513<=SI513;
out514<=SI514;
out515<=SI515;
out516<=SI516;
out517<=SI517;
out518<=SI518;
out519<=SI519;
out520<=SI520;
out521<=SI521;
out522<=SI522;
out523<=SI523;
out524<=SI524;
out525<=SI525;
out526<=SI526;
out527<=SI527;
out528<=SI528;
out529<=SI529;
out530<=SI530;
out531<=SI531;
out532<=SI532;
out533<=SI533;
out534<=SI534;
out535<=SI535;
out536<=SI536;
out537<=SI537;
out538<=SI538;
out539<=SI539;
out540<=SI540;
out541<=SI541;
out542<=SI542;
out543<=SI543;
out544<=SI544;
out545<=SI545;
out546<=SI546;
out547<=SI547;
out548<=SI548;
out549<=SI549;
out550<=SI550;
out551<=SI551;
out552<=SI552;
out553<=SI553;
out554<=SI554;
out555<=SI555;
out556<=SI556;
out557<=SI557;
out558<=SI558;
out559<=SI559;
out560<=SI560;
out561<=SI561;
out562<=SI562;
out563<=SI563;
out564<=SI564;
out565<=SI565;
out566<=SI566;
out567<=SI567;
out568<=SI568;
out569<=SI569;
out570<=SI570;
out571<=SI571;
out572<=SI572;
out573<=SI573;
out574<=SI574;
out575<=SI575;
out576<=SI576;
out577<=SI577;
out578<=SI578;
out579<=SI579;
out580<=SI580;
out581<=SI581;
out582<=SI582;
out583<=SI583;
out584<=SI584;
out585<=SI585;
out586<=SI586;
out587<=SI587;
out588<=SI588;
out589<=SI589;
out590<=SI590;
out591<=SI591;
out592<=SI592;
out593<=SI593;
out594<=SI594;
out595<=SI595;
out596<=SI596;
out597<=SI597;
out598<=SI598;
out599<=SI599;
out600<=SI600;
out601<=SI601;
out602<=SI602;
out603<=SI603;
out604<=SI604;
out605<=SI605;
out606<=SI606;
out607<=SI607;
out608<=SI608;
out609<=SI609;
out610<=SI610;
out611<=SI611;
out612<=SI612;
out613<=SI613;
out614<=SI614;
out615<=SI615;
out616<=SI616;
out617<=SI617;
out618<=SI618;
out619<=SI619;
out620<=SI620;
out621<=SI621;
out622<=SI622;
out623<=SI623;
out624<=SI624;
out625<=SI625;
out626<=SI626;
out627<=SI627;
out628<=SI628;
out629<=SI629;
out630<=SI630;
out631<=SI631;
out632<=SI632;
out633<=SI633;
out634<=SI634;
out635<=SI635;
out636<=SI636;
out637<=SI637;
out638<=SI638;
out639<=SI639;
out640<=SI640;
out641<=SI641;
out642<=SI642;
out643<=SI643;
out644<=SI644;
out645<=SI645;
out646<=SI646;
out647<=SI647;
out648<=SI648;
out649<=SI649;
out650<=SI650;
out651<=SI651;
out652<=SI652;
out653<=SI653;
out654<=SI654;
out655<=SI655;
out656<=SI656;
out657<=SI657;
out658<=SI658;
out659<=SI659;
out660<=SI660;
out661<=SI661;
out662<=SI662;
out663<=SI663;
out664<=SI664;
out665<=SI665;
out666<=SI666;
out667<=SI667;
out668<=SI668;
out669<=SI669;
out670<=SI670;
out671<=SI671;
out672<=SI672;
out673<=SI673;
out674<=SI674;
out675<=SI675;
out676<=SI676;
out677<=SI677;
out678<=SI678;
out679<=SI679;
out680<=SI680;
out681<=SI681;
out682<=SI682;
out683<=SI683;
out684<=SI684;
out685<=SI685;
out686<=SI686;
out687<=SI687;
out688<=SI688;
out689<=SI689;
out690<=SI690;
out691<=SI691;
out692<=SI692;
out693<=SI693;
out694<=SI694;
out695<=SI695;
out696<=SI696;
out697<=SI697;
out698<=SI698;
out699<=SI699;
out700<=SI700;
out701<=SI701;
out702<=SI702;
out703<=SI703;
out704<=SI704;
out705<=SI705;
out706<=SI706;
out707<=SI707;
out708<=SI708;
out709<=SI709;
out710<=SI710;
out711<=SI711;
out712<=SI712;
out713<=SI713;
out714<=SI714;
out715<=SI715;
out716<=SI716;
out717<=SI717;
out718<=SI718;
out719<=SI719;
out720<=SI720;
out721<=SI721;
out722<=SI722;
out723<=SI723;
out724<=SI724;
out725<=SI725;
out726<=SI726;
out727<=SI727;
out728<=SI728;
out729<=SI729;
out730<=SI730;
out731<=SI731;
out732<=SI732;
out733<=SI733;
out734<=SI734;
out735<=SI735;
out736<=SI736;
out737<=SI737;
out738<=SI738;
out739<=SI739;
out740<=SI740;
out741<=SI741;
out742<=SI742;
out743<=SI743;
out744<=SI744;
out745<=SI745;
out746<=SI746;
out747<=SI747;
out748<=SI748;
out749<=SI749;
out750<=SI750;
out751<=SI751;
out752<=SI752;
out753<=SI753;
out754<=SI754;
out755<=SI755;
out756<=SI756;
out757<=SI757;
out758<=SI758;
out759<=SI759;
out760<=SI760;
out761<=SI761;
out762<=SI762;
out763<=SI763;
out764<=SI764;
out765<=SI765;
out766<=SI766;
out767<=SI767;
out768<=SI768;
out769<=SI769;
out770<=SI770;
out771<=SI771;
out772<=SI772;
out773<=SI773;
out774<=SI774;
out775<=SI775;
out776<=SI776;
out777<=SI777;
out778<=SI778;
out779<=SI779;
out780<=SI780;
out781<=SI781;
out782<=SI782;
out783<=SI783;
out784<=SI784;
out785<=SI785;
out786<=SI786;
out787<=SI787;
out788<=SI788;
out789<=SI789;
out790<=SI790;
out791<=SI791;
out792<=SI792;
out793<=SI793;
out794<=SI794;
out795<=SI795;
out796<=SI796;
out797<=SI797;
out798<=SI798;
out799<=SI799;
out800<=SI800;
out801<=SI801;
out802<=SI802;
out803<=SI803;
out804<=SI804;
out805<=SI805;
out806<=SI806;
out807<=SI807;
out808<=SI808;
out809<=SI809;
out810<=SI810;
out811<=SI811;
out812<=SI812;
out813<=SI813;
out814<=SI814;
out815<=SI815;
out816<=SI816;
out817<=SI817;
out818<=SI818;
out819<=SI819;
out820<=SI820;
out821<=SI821;
out822<=SI822;
out823<=SI823;
out824<=SI824;
out825<=SI825;
out826<=SI826;
out827<=SI827;
out828<=SI828;
out829<=SI829;
out830<=SI830;
out831<=SI831;
out832<=SI832;
out833<=SI833;
out834<=SI834;
out835<=SI835;
out836<=SI836;
out837<=SI837;
out838<=SI838;
out839<=SI839;
out840<=SI840;
out841<=SI841;
out842<=SI842;
out843<=SI843;
out844<=SI844;
out845<=SI845;
out846<=SI846;
out847<=SI847;
out848<=SI848;
out849<=SI849;
out850<=SI850;
out851<=SI851;
out852<=SI852;
out853<=SI853;
out854<=SI854;
out855<=SI855;
out856<=SI856;
out857<=SI857;
out858<=SI858;
out859<=SI859;
out860<=SI860;
out861<=SI861;
out862<=SI862;
out863<=SI863;
out864<=SI864;
out865<=SI865;
out866<=SI866;
out867<=SI867;
out868<=SI868;
out869<=SI869;
out870<=SI870;
out871<=SI871;
out872<=SI872;
out873<=SI873;
out874<=SI874;
out875<=SI875;
out876<=SI876;
out877<=SI877;
out878<=SI878;
out879<=SI879;
out880<=SI880;
out881<=SI881;
out882<=SI882;
out883<=SI883;
out884<=SI884;
out885<=SI885;
out886<=SI886;
out887<=SI887;
out888<=SI888;
out889<=SI889;
out890<=SI890;
out891<=SI891;
out892<=SI892;
out893<=SI893;
out894<=SI894;
out895<=SI895;
out896<=SI896;
out897<=SI897;
out898<=SI898;
out899<=SI899;
out900<=SI900;
out901<=SI901;
out902<=SI902;
out903<=SI903;
out904<=SI904;
out905<=SI905;
out906<=SI906;
out907<=SI907;
out908<=SI908;
out909<=SI909;
out910<=SI910;
out911<=SI911;
out912<=SI912;
out913<=SI913;
out914<=SI914;
out915<=SI915;
out916<=SI916;
out917<=SI917;
out918<=SI918;
out919<=SI919;
out920<=SI920;
out921<=SI921;
out922<=SI922;
out923<=SI923;
out924<=SI924;
out925<=SI925;
out926<=SI926;
out927<=SI927;
out928<=SI928;
out929<=SI929;
out930<=SI930;
out931<=SI931;
out932<=SI932;
out933<=SI933;
out934<=SI934;
out935<=SI935;
out936<=SI936;
out937<=SI937;
out938<=SI938;
out939<=SI939;
out940<=SI940;
out941<=SI941;
out942<=SI942;
out943<=SI943;
out944<=SI944;
out945<=SI945;
out946<=SI946;
out947<=SI947;
out948<=SI948;
out949<=SI949;
out950<=SI950;
out951<=SI951;
out952<=SI952;
out953<=SI953;
out954<=SI954;
out955<=SI955;
out956<=SI956;
out957<=SI957;
out958<=SI958;
out959<=SI959;
out960<=SI960;
out961<=SI961;
out962<=SI962;
out963<=SI963;
out964<=SI964;
out965<=SI965;
out966<=SI966;
out967<=SI967;
out968<=SI968;
out969<=SI969;
out970<=SI970;
out971<=SI971;
out972<=SI972;
out973<=SI973;
out974<=SI974;
out975<=SI975;
out976<=SI976;
out977<=SI977;
out978<=SI978;
out979<=SI979;
out980<=SI980;
out981<=SI981;
out982<=SI982;
out983<=SI983;
out984<=SI984;
out985<=SI985;
out986<=SI986;
out987<=SI987;
out988<=SI988;
out989<=SI989;
out990<=SI990;
out991<=SI991;
out992<=SI992;
out993<=SI993;
out994<=SI994;
out995<=SI995;
out996<=SI996;
out997<=SI997;
out998<=SI998;
out999<=SI999;
out1000<=SI1000;
out1001<=SI1001;
out1002<=SI1002;
out1003<=SI1003;
out1004<=SI1004;
out1005<=SI1005;
out1006<=SI1006;
out1007<=SI1007;
out1008<=SI1008;
out1009<=SI1009;
out1010<=SI1010;
out1011<=SI1011;
out1012<=SI1012;
out1013<=SI1013;
out1014<=SI1014;
out1015<=SI1015;
out1016<=SI1016;
out1017<=SI1017;
out1018<=SI1018;
out1019<=SI1019;
out1020<=SI1020;
out1021<=SI1021;
out1022<=SI1022;
out1023<=SI1023;
out1024<=SI1024;
out1025<=SI1025;
out1026<=SI1026;
out1027<=SI1027;
out1028<=SI1028;
out1029<=SI1029;
out1030<=SI1030;
out1031<=SI1031;
out1032<=SI1032;
out1033<=SI1033;
out1034<=SI1034;
out1035<=SI1035;
out1036<=SI1036;
out1037<=SI1037;
out1038<=SI1038;
out1039<=SI1039;
out1040<=SI1040;
out1041<=SI1041;
out1042<=SI1042;
out1043<=SI1043;
out1044<=SI1044;
out1045<=SI1045;
out1046<=SI1046;
out1047<=SI1047;
out1048<=SI1048;
out1049<=SI1049;
out1050<=SI1050;
out1051<=SI1051;
out1052<=SI1052;
out1053<=SI1053;
out1054<=SI1054;
out1055<=SI1055;
out1056<=SI1056;
out1057<=SI1057;
out1058<=SI1058;
out1059<=SI1059;
out1060<=SI1060;
out1061<=SI1061;
out1062<=SI1062;
out1063<=SI1063;
out1064<=SI1064;
out1065<=SI1065;
out1066<=SI1066;
out1067<=SI1067;
out1068<=SI1068;
out1069<=SI1069;
out1070<=SI1070;
out1071<=SI1071;
out1072<=SI1072;
out1073<=SI1073;
out1074<=SI1074;
out1075<=SI1075;
out1076<=SI1076;
out1077<=SI1077;
out1078<=SI1078;
out1079<=SI1079;
out1080<=SI1080;
out1081<=SI1081;
out1082<=SI1082;
out1083<=SI1083;
out1084<=SI1084;
out1085<=SI1085;
out1086<=SI1086;
out1087<=SI1087;
out1088<=SI1088;
out1089<=SI1089;
out1090<=SI1090;
out1091<=SI1091;
out1092<=SI1092;
out1093<=SI1093;
out1094<=SI1094;
out1095<=SI1095;
out1096<=SI1096;
out1097<=SI1097;
out1098<=SI1098;
out1099<=SI1099;
out1100<=SI1100;
out1101<=SI1101;
out1102<=SI1102;
out1103<=SI1103;
out1104<=SI1104;
out1105<=SI1105;
out1106<=SI1106;
out1107<=SI1107;
out1108<=SI1108;
out1109<=SI1109;
out1110<=SI1110;
out1111<=SI1111;
out1112<=SI1112;
out1113<=SI1113;
out1114<=SI1114;
out1115<=SI1115;
out1116<=SI1116;
out1117<=SI1117;
out1118<=SI1118;
out1119<=SI1119;
out1120<=SI1120;
out1121<=SI1121;
out1122<=SI1122;
out1123<=SI1123;
out1124<=SI1124;
out1125<=SI1125;
out1126<=SI1126;
out1127<=SI1127;
out1128<=SI1128;
out1129<=SI1129;
out1130<=SI1130;
out1131<=SI1131;
out1132<=SI1132;
out1133<=SI1133;
out1134<=SI1134;
out1135<=SI1135;
out1136<=SI1136;
out1137<=SI1137;
out1138<=SI1138;
out1139<=SI1139;
out1140<=SI1140;
out1141<=SI1141;
out1142<=SI1142;
out1143<=SI1143;
out1144<=SI1144;
out1145<=SI1145;
out1146<=SI1146;
out1147<=SI1147;
out1148<=SI1148;
out1149<=SI1149;
out1150<=SI1150;
out1151<=SI1151;
out1152<=SI1152;
out1153<=SI1153;
out1154<=SI1154;
out1155<=SI1155;
out1156<=SI1156;
out1157<=SI1157;
out1158<=SI1158;
out1159<=SI1159;
out1160<=SI1160;
out1161<=SI1161;
out1162<=SI1162;
out1163<=SI1163;
out1164<=SI1164;
out1165<=SI1165;
out1166<=SI1166;
out1167<=SI1167;
out1168<=SI1168;
out1169<=SI1169;
out1170<=SI1170;
out1171<=SI1171;
out1172<=SI1172;
out1173<=SI1173;
out1174<=SI1174;
out1175<=SI1175;
out1176<=SI1176;
out1177<=SI1177;
out1178<=SI1178;
out1179<=SI1179;
out1180<=SI1180;
out1181<=SI1181;
out1182<=SI1182;
out1183<=SI1183;
out1184<=SI1184;
out1185<=SI1185;
out1186<=SI1186;
out1187<=SI1187;
out1188<=SI1188;
out1189<=SI1189;
out1190<=SI1190;
out1191<=SI1191;
out1192<=SI1192;
out1193<=SI1193;
out1194<=SI1194;
out1195<=SI1195;
out1196<=SI1196;
out1197<=SI1197;
out1198<=SI1198;
out1199<=SI1199;
out1200<=SI1200;
out1201<=SI1201;
out1202<=SI1202;
out1203<=SI1203;
out1204<=SI1204;
out1205<=SI1205;
out1206<=SI1206;
out1207<=SI1207;
out1208<=SI1208;
out1209<=SI1209;
out1210<=SI1210;
out1211<=SI1211;
out1212<=SI1212;
out1213<=SI1213;
out1214<=SI1214;
out1215<=SI1215;
out1216<=SI1216;
out1217<=SI1217;
out1218<=SI1218;
out1219<=SI1219;
out1220<=SI1220;
out1221<=SI1221;
out1222<=SI1222;
out1223<=SI1223;
out1224<=SI1224;
out1225<=SI1225;
out1226<=SI1226;
out1227<=SI1227;
out1228<=SI1228;
out1229<=SI1229;
out1230<=SI1230;
out1231<=SI1231;
out1232<=SI1232;
out1233<=SI1233;
out1234<=SI1234;
out1235<=SI1235;
out1236<=SI1236;
out1237<=SI1237;
out1238<=SI1238;
out1239<=SI1239;
out1240<=SI1240;
out1241<=SI1241;
out1242<=SI1242;
out1243<=SI1243;
out1244<=SI1244;
out1245<=SI1245;
out1246<=SI1246;
out1247<=SI1247;
out1248<=SI1248;
out1249<=SI1249;
out1250<=SI1250;
out1251<=SI1251;
out1252<=SI1252;
out1253<=SI1253;
out1254<=SI1254;
out1255<=SI1255;
out1256<=SI1256;
out1257<=SI1257;
out1258<=SI1258;
out1259<=SI1259;
out1260<=SI1260;
out1261<=SI1261;
out1262<=SI1262;
out1263<=SI1263;
out1264<=SI1264;
out1265<=SI1265;
out1266<=SI1266;
out1267<=SI1267;
out1268<=SI1268;
out1269<=SI1269;
out1270<=SI1270;
out1271<=SI1271;
out1272<=SI1272;
out1273<=SI1273;
out1274<=SI1274;
out1275<=SI1275;
out1276<=SI1276;
out1277<=SI1277;
out1278<=SI1278;
out1279<=SI1279;
out1280<=SI1280;
out1281<=SI1281;
out1282<=SI1282;
out1283<=SI1283;
out1284<=SI1284;
out1285<=SI1285;
out1286<=SI1286;
out1287<=SI1287;
out1288<=SI1288;
out1289<=SI1289;
out1290<=SI1290;
out1291<=SI1291;
out1292<=SI1292;
out1293<=SI1293;
out1294<=SI1294;
out1295<=SI1295;
out1296<=SI1296;
out1297<=SI1297;
out1298<=SI1298;
out1299<=SI1299;
out1300<=SI1300;
out1301<=SI1301;
out1302<=SI1302;
out1303<=SI1303;
out1304<=SI1304;
out1305<=SI1305;
out1306<=SI1306;
out1307<=SI1307;
out1308<=SI1308;
out1309<=SI1309;
out1310<=SI1310;
out1311<=SI1311;
out1312<=SI1312;
out1313<=SI1313;
out1314<=SI1314;
out1315<=SI1315;
out1316<=SI1316;
out1317<=SI1317;
out1318<=SI1318;
out1319<=SI1319;
out1320<=SI1320;
out1321<=SI1321;
out1322<=SI1322;
out1323<=SI1323;
out1324<=SI1324;
out1325<=SI1325;
out1326<=SI1326;
out1327<=SI1327;
out1328<=SI1328;
out1329<=SI1329;
out1330<=SI1330;
out1331<=SI1331;
out1332<=SI1332;
out1333<=SI1333;
out1334<=SI1334;
out1335<=SI1335;
out1336<=SI1336;
out1337<=SI1337;
out1338<=SI1338;
out1339<=SI1339;
out1340<=SI1340;
out1341<=SI1341;
out1342<=SI1342;
out1343<=SI1343;
out1344<=SI1344;
out1345<=SI1345;
out1346<=SI1346;
out1347<=SI1347;
out1348<=SI1348;
out1349<=SI1349;
out1350<=SI1350;
out1351<=SI1351;
out1352<=SI1352;
out1353<=SI1353;
out1354<=SI1354;
out1355<=SI1355;
out1356<=SI1356;
out1357<=SI1357;
out1358<=SI1358;
out1359<=SI1359;
out1360<=SI1360;
out1361<=SI1361;
out1362<=SI1362;
out1363<=SI1363;
out1364<=SI1364;
out1365<=SI1365;
out1366<=SI1366;
out1367<=SI1367;
out1368<=SI1368;
out1369<=SI1369;
out1370<=SI1370;
out1371<=SI1371;
out1372<=SI1372;
out1373<=SI1373;
out1374<=SI1374;
out1375<=SI1375;
out1376<=SI1376;
out1377<=SI1377;
out1378<=SI1378;
out1379<=SI1379;
out1380<=SI1380;
out1381<=SI1381;
out1382<=SI1382;
out1383<=SI1383;
out1384<=SI1384;
out1385<=SI1385;
out1386<=SI1386;
out1387<=SI1387;
out1388<=SI1388;
out1389<=SI1389;
out1390<=SI1390;
out1391<=SI1391;
out1392<=SI1392;
out1393<=SI1393;
out1394<=SI1394;
out1395<=SI1395;
out1396<=SI1396;
out1397<=SI1397;
out1398<=SI1398;
out1399<=SI1399;
out1400<=SI1400;
out1401<=SI1401;
out1402<=SI1402;
out1403<=SI1403;
out1404<=SI1404;
out1405<=SI1405;
out1406<=SI1406;
out1407<=SI1407;
out1408<=SI1408;
out1409<=SI1409;
out1410<=SI1410;
out1411<=SI1411;
out1412<=SI1412;
out1413<=SI1413;
out1414<=SI1414;
out1415<=SI1415;
out1416<=SI1416;
out1417<=SI1417;
out1418<=SI1418;
out1419<=SI1419;
out1420<=SI1420;
out1421<=SI1421;
out1422<=SI1422;
out1423<=SI1423;
out1424<=SI1424;
out1425<=SI1425;
out1426<=SI1426;
out1427<=SI1427;
out1428<=SI1428;
out1429<=SI1429;
out1430<=SI1430;
out1431<=SI1431;
out1432<=SI1432;
out1433<=SI1433;
out1434<=SI1434;
out1435<=SI1435;
out1436<=SI1436;
out1437<=SI1437;
out1438<=SI1438;
out1439<=SI1439;
out1440<=SI1440;
out1441<=SI1441;
out1442<=SI1442;
out1443<=SI1443;
out1444<=SI1444;
out1445<=SI1445;
out1446<=SI1446;
out1447<=SI1447;
out1448<=SI1448;
out1449<=SI1449;
out1450<=SI1450;
out1451<=SI1451;
out1452<=SI1452;
out1453<=SI1453;
out1454<=SI1454;
out1455<=SI1455;
out1456<=SI1456;
out1457<=SI1457;
out1458<=SI1458;
out1459<=SI1459;
out1460<=SI1460;
out1461<=SI1461;
out1462<=SI1462;
out1463<=SI1463;
out1464<=SI1464;
out1465<=SI1465;
out1466<=SI1466;
out1467<=SI1467;
out1468<=SI1468;
out1469<=SI1469;
out1470<=SI1470;
out1471<=SI1471;
out1472<=SI1472;
out1473<=SI1473;
out1474<=SI1474;
out1475<=SI1475;
out1476<=SI1476;
out1477<=SI1477;
out1478<=SI1478;
out1479<=SI1479;
out1480<=SI1480;
out1481<=SI1481;
out1482<=SI1482;
out1483<=SI1483;
out1484<=SI1484;
out1485<=SI1485;
out1486<=SI1486;
out1487<=SI1487;
out1488<=SI1488;
out1489<=SI1489;
out1490<=SI1490;
out1491<=SI1491;
out1492<=SI1492;
out1493<=SI1493;
out1494<=SI1494;
out1495<=SI1495;
out1496<=SI1496;
out1497<=SI1497;
out1498<=SI1498;
out1499<=SI1499;
out1500<=SI1500;
out1501<=SI1501;
out1502<=SI1502;
out1503<=SI1503;
out1504<=SI1504;
out1505<=SI1505;
out1506<=SI1506;
out1507<=SI1507;
out1508<=SI1508;
out1509<=SI1509;
out1510<=SI1510;
out1511<=SI1511;
out1512<=SI1512;
out1513<=SI1513;
out1514<=SI1514;
out1515<=SI1515;
out1516<=SI1516;
out1517<=SI1517;
out1518<=SI1518;
out1519<=SI1519;
out1520<=SI1520;
out1521<=SI1521;
out1522<=SI1522;
out1523<=SI1523;
out1524<=SI1524;
out1525<=SI1525;
out1526<=SI1526;
out1527<=SI1527;
out1528<=SI1528;
out1529<=SI1529;
out1530<=SI1530;
out1531<=SI1531;
out1532<=SI1532;
out1533<=SI1533;
out1534<=SI1534;
out1535<=SI1535;
out1536<=SI1536;
out1537<=SI1537;
out1538<=SI1538;
out1539<=SI1539;
out1540<=SI1540;
out1541<=SI1541;
out1542<=SI1542;
out1543<=SI1543;
out1544<=SI1544;
out1545<=SI1545;
out1546<=SI1546;
out1547<=SI1547;
out1548<=SI1548;
out1549<=SI1549;
out1550<=SI1550;
out1551<=SI1551;
out1552<=SI1552;
out1553<=SI1553;
out1554<=SI1554;
out1555<=SI1555;
out1556<=SI1556;
out1557<=SI1557;
out1558<=SI1558;
out1559<=SI1559;
out1560<=SI1560;
out1561<=SI1561;
out1562<=SI1562;
out1563<=SI1563;
out1564<=SI1564;
out1565<=SI1565;
out1566<=SI1566;
out1567<=SI1567;
out1568<=SI1568;
out1569<=SI1569;
out1570<=SI1570;
out1571<=SI1571;
out1572<=SI1572;
out1573<=SI1573;
out1574<=SI1574;
out1575<=SI1575;
out1576<=SI1576;
out1577<=SI1577;
out1578<=SI1578;
out1579<=SI1579;
out1580<=SI1580;
out1581<=SI1581;
out1582<=SI1582;
out1583<=SI1583;
out1584<=SI1584;
out1585<=SI1585;
out1586<=SI1586;
out1587<=SI1587;
out1588<=SI1588;
out1589<=SI1589;
out1590<=SI1590;
out1591<=SI1591;
out1592<=SI1592;
out1593<=SI1593;
out1594<=SI1594;
out1595<=SI1595;
out1596<=SI1596;
out1597<=SI1597;
out1598<=SI1598;
out1599<=SI1599;
out1600<=SI1600;
out1601<=SI1601;
out1602<=SI1602;
out1603<=SI1603;
out1604<=SI1604;
out1605<=SI1605;
out1606<=SI1606;
out1607<=SI1607;
out1608<=SI1608;
out1609<=SI1609;
out1610<=SI1610;
out1611<=SI1611;
out1612<=SI1612;
out1613<=SI1613;
out1614<=SI1614;
out1615<=SI1615;
out1616<=SI1616;
out1617<=SI1617;
out1618<=SI1618;
out1619<=SI1619;
out1620<=SI1620;
out1621<=SI1621;
out1622<=SI1622;
out1623<=SI1623;
out1624<=SI1624;
out1625<=SI1625;
out1626<=SI1626;
out1627<=SI1627;
out1628<=SI1628;
out1629<=SI1629;
out1630<=SI1630;
out1631<=SI1631;
out1632<=SI1632;
out1633<=SI1633;
out1634<=SI1634;
out1635<=SI1635;
out1636<=SI1636;
out1637<=SI1637;
out1638<=SI1638;
out1639<=SI1639;
out1640<=SI1640;
out1641<=SI1641;
out1642<=SI1642;
out1643<=SI1643;
out1644<=SI1644;
out1645<=SI1645;
out1646<=SI1646;
out1647<=SI1647;
out1648<=SI1648;
out1649<=SI1649;
out1650<=SI1650;
out1651<=SI1651;
out1652<=SI1652;
out1653<=SI1653;
out1654<=SI1654;
out1655<=SI1655;
out1656<=SI1656;
out1657<=SI1657;
out1658<=SI1658;
out1659<=SI1659;
out1660<=SI1660;
out1661<=SI1661;
out1662<=SI1662;
out1663<=SI1663;
out1664<=SI1664;
out1665<=SI1665;
out1666<=SI1666;
out1667<=SI1667;
out1668<=SI1668;
out1669<=SI1669;
out1670<=SI1670;
out1671<=SI1671;
out1672<=SI1672;
out1673<=SI1673;
out1674<=SI1674;
out1675<=SI1675;
out1676<=SI1676;
out1677<=SI1677;
out1678<=SI1678;
out1679<=SI1679;
out1680<=SI1680;
out1681<=SI1681;
out1682<=SI1682;
out1683<=SI1683;
out1684<=SI1684;
out1685<=SI1685;
out1686<=SI1686;
out1687<=SI1687;
out1688<=SI1688;
out1689<=SI1689;
out1690<=SI1690;
out1691<=SI1691;
out1692<=SI1692;
out1693<=SI1693;
out1694<=SI1694;
out1695<=SI1695;
out1696<=SI1696;
out1697<=SI1697;
out1698<=SI1698;
out1699<=SI1699;
out1700<=SI1700;
out1701<=SI1701;
out1702<=SI1702;
out1703<=SI1703;
out1704<=SI1704;
out1705<=SI1705;
out1706<=SI1706;
out1707<=SI1707;
out1708<=SI1708;
out1709<=SI1709;
out1710<=SI1710;
out1711<=SI1711;
out1712<=SI1712;
out1713<=SI1713;
out1714<=SI1714;
out1715<=SI1715;
out1716<=SI1716;
out1717<=SI1717;
out1718<=SI1718;
out1719<=SI1719;
out1720<=SI1720;
out1721<=SI1721;
out1722<=SI1722;
out1723<=SI1723;
out1724<=SI1724;
out1725<=SI1725;
out1726<=SI1726;
out1727<=SI1727;
out1728<=SI1728;
out1729<=SI1729;
out1730<=SI1730;
out1731<=SI1731;
out1732<=SI1732;
out1733<=SI1733;
out1734<=SI1734;
out1735<=SI1735;
out1736<=SI1736;
out1737<=SI1737;
out1738<=SI1738;
out1739<=SI1739;
out1740<=SI1740;
out1741<=SI1741;
out1742<=SI1742;
out1743<=SI1743;
out1744<=SI1744;
out1745<=SI1745;
out1746<=SI1746;
out1747<=SI1747;
out1748<=SI1748;
out1749<=SI1749;
out1750<=SI1750;
out1751<=SI1751;
out1752<=SI1752;
out1753<=SI1753;
out1754<=SI1754;
out1755<=SI1755;
out1756<=SI1756;
out1757<=SI1757;
out1758<=SI1758;
out1759<=SI1759;
out1760<=SI1760;
out1761<=SI1761;
out1762<=SI1762;
out1763<=SI1763;
out1764<=SI1764;
out1765<=SI1765;
out1766<=SI1766;
out1767<=SI1767;
out1768<=SI1768;
out1769<=SI1769;
out1770<=SI1770;
out1771<=SI1771;
out1772<=SI1772;
out1773<=SI1773;
out1774<=SI1774;
out1775<=SI1775;
out1776<=SI1776;
out1777<=SI1777;
out1778<=SI1778;
out1779<=SI1779;
out1780<=SI1780;
out1781<=SI1781;
out1782<=SI1782;
out1783<=SI1783;
out1784<=SI1784;
out1785<=SI1785;
out1786<=SI1786;
out1787<=SI1787;
out1788<=SI1788;
out1789<=SI1789;
out1790<=SI1790;
out1791<=SI1791;
out1792<=SI1792;
out1793<=SI1793;
out1794<=SI1794;
out1795<=SI1795;
out1796<=SI1796;
out1797<=SI1797;
out1798<=SI1798;
out1799<=SI1799;
out1800<=SI1800;
out1801<=SI1801;
out1802<=SI1802;
out1803<=SI1803;
out1804<=SI1804;
out1805<=SI1805;
out1806<=SI1806;
out1807<=SI1807;
out1808<=SI1808;
out1809<=SI1809;
out1810<=SI1810;
out1811<=SI1811;
out1812<=SI1812;
out1813<=SI1813;
out1814<=SI1814;
out1815<=SI1815;
out1816<=SI1816;
out1817<=SI1817;
out1818<=SI1818;
out1819<=SI1819;
out1820<=SI1820;
out1821<=SI1821;
out1822<=SI1822;
out1823<=SI1823;
out1824<=SI1824;
out1825<=SI1825;
out1826<=SI1826;
out1827<=SI1827;
out1828<=SI1828;
out1829<=SI1829;
out1830<=SI1830;
out1831<=SI1831;
out1832<=SI1832;
out1833<=SI1833;
out1834<=SI1834;
out1835<=SI1835;
out1836<=SI1836;
out1837<=SI1837;
out1838<=SI1838;
out1839<=SI1839;
out1840<=SI1840;
out1841<=SI1841;
out1842<=SI1842;
out1843<=SI1843;
out1844<=SI1844;
out1845<=SI1845;
out1846<=SI1846;
out1847<=SI1847;
out1848<=SI1848;
out1849<=SI1849;
out1850<=SI1850;
out1851<=SI1851;
out1852<=SI1852;
out1853<=SI1853;
out1854<=SI1854;
out1855<=SI1855;
out1856<=SI1856;
out1857<=SI1857;
out1858<=SI1858;
out1859<=SI1859;
out1860<=SI1860;
out1861<=SI1861;
out1862<=SI1862;
out1863<=SI1863;
out1864<=SI1864;
out1865<=SI1865;
out1866<=SI1866;
out1867<=SI1867;
out1868<=SI1868;
out1869<=SI1869;
out1870<=SI1870;
out1871<=SI1871;
out1872<=SI1872;
out1873<=SI1873;
out1874<=SI1874;
out1875<=SI1875;
out1876<=SI1876;
out1877<=SI1877;
out1878<=SI1878;
out1879<=SI1879;
out1880<=SI1880;
out1881<=SI1881;
out1882<=SI1882;
out1883<=SI1883;
out1884<=SI1884;
out1885<=SI1885;
out1886<=SI1886;
out1887<=SI1887;
out1888<=SI1888;
out1889<=SI1889;
out1890<=SI1890;
out1891<=SI1891;
out1892<=SI1892;
out1893<=SI1893;
out1894<=SI1894;
out1895<=SI1895;
out1896<=SI1896;
out1897<=SI1897;
out1898<=SI1898;
out1899<=SI1899;
out1900<=SI1900;
out1901<=SI1901;
out1902<=SI1902;
out1903<=SI1903;
out1904<=SI1904;
out1905<=SI1905;
out1906<=SI1906;
out1907<=SI1907;
out1908<=SI1908;
out1909<=SI1909;
out1910<=SI1910;
out1911<=SI1911;
out1912<=SI1912;
out1913<=SI1913;
out1914<=SI1914;
out1915<=SI1915;
out1916<=SI1916;
out1917<=SI1917;
out1918<=SI1918;
out1919<=SI1919;
out1920<=SI1920;
out1921<=SI1921;
out1922<=SI1922;
out1923<=SI1923;
out1924<=SI1924;
out1925<=SI1925;
out1926<=SI1926;
out1927<=SI1927;
out1928<=SI1928;
out1929<=SI1929;
out1930<=SI1930;
out1931<=SI1931;
out1932<=SI1932;
out1933<=SI1933;
out1934<=SI1934;
out1935<=SI1935;
out1936<=SI1936;
out1937<=SI1937;
out1938<=SI1938;
out1939<=SI1939;
out1940<=SI1940;
out1941<=SI1941;
out1942<=SI1942;
out1943<=SI1943;
out1944<=SI1944;
out1945<=SI1945;
out1946<=SI1946;
out1947<=SI1947;
out1948<=SI1948;
out1949<=SI1949;
out1950<=SI1950;
out1951<=SI1951;
out1952<=SI1952;
out1953<=SI1953;
out1954<=SI1954;
out1955<=SI1955;
out1956<=SI1956;
out1957<=SI1957;
out1958<=SI1958;
out1959<=SI1959;
out1960<=SI1960;
out1961<=SI1961;
out1962<=SI1962;
out1963<=SI1963;
out1964<=SI1964;
out1965<=SI1965;
out1966<=SI1966;
out1967<=SI1967;
out1968<=SI1968;
out1969<=SI1969;
out1970<=SI1970;
out1971<=SI1971;
out1972<=SI1972;
out1973<=SI1973;
out1974<=SI1974;
out1975<=SI1975;
out1976<=SI1976;
out1977<=SI1977;
out1978<=SI1978;
out1979<=SI1979;
out1980<=SI1980;
out1981<=SI1981;
out1982<=SI1982;
out1983<=SI1983;
out1984<=SI1984;
out1985<=SI1985;
out1986<=SI1986;
out1987<=SI1987;
out1988<=SI1988;
out1989<=SI1989;
out1990<=SI1990;
out1991<=SI1991;
out1992<=SI1992;
out1993<=SI1993;
out1994<=SI1994;
out1995<=SI1995;
out1996<=SI1996;
out1997<=SI1997;
out1998<=SI1998;
out1999<=SI1999;
out2000<=SI2000;
out2001<=SI2001;
out2002<=SI2002;
out2003<=SI2003;
out2004<=SI2004;
out2005<=SI2005;
out2006<=SI2006;
out2007<=SI2007;
out2008<=SI2008;
out2009<=SI2009;
out2010<=SI2010;
out2011<=SI2011;
out2012<=SI2012;
out2013<=SI2013;
out2014<=SI2014;
out2015<=SI2015;
out2016<=SI2016;
out2017<=SI2017;
out2018<=SI2018;
out2019<=SI2019;
out2020<=SI2020;
out2021<=SI2021;
out2022<=SI2022;
out2023<=SI2023;
out2024<=SI2024;
out2025<=SI2025;
out2026<=SI2026;
out2027<=SI2027;
out2028<=SI2028;
out2029<=SI2029;
out2030<=SI2030;
out2031<=SI2031;
out2032<=SI2032;
out2033<=SI2033;
out2034<=SI2034;
out2035<=SI2035;
out2036<=SI2036;
out2037<=SI2037;
out2038<=SI2038;
out2039<=SI2039;
out2040<=SI2040;
out2041<=SI2041;
out2042<=SI2042;
out2043<=SI2043;
out2044<=SI2044;
out2045<=SI2045;
out2046<=SI2046;
out2047<=SI2047;
out2048<=SI2048;
out2049<=SI2049;
out2050<=SI2050;
out2051<=SI2051;
out2052<=SI2052;
out2053<=SI2053;
out2054<=SI2054;
out2055<=SI2055;
out2056<=SI2056;
out2057<=SI2057;
out2058<=SI2058;
out2059<=SI2059;
out2060<=SI2060;
out2061<=SI2061;
out2062<=SI2062;
out2063<=SI2063;
out2064<=SI2064;
out2065<=SI2065;
out2066<=SI2066;
out2067<=SI2067;
out2068<=SI2068;
out2069<=SI2069;
out2070<=SI2070;
out2071<=SI2071;
out2072<=SI2072;
out2073<=SI2073;
out2074<=SI2074;
out2075<=SI2075;
out2076<=SI2076;
out2077<=SI2077;
out2078<=SI2078;
out2079<=SI2079;
out2080<=SI2080;
out2081<=SI2081;
out2082<=SI2082;
out2083<=SI2083;
out2084<=SI2084;
out2085<=SI2085;
out2086<=SI2086;
out2087<=SI2087;
out2088<=SI2088;
out2089<=SI2089;
out2090<=SI2090;
out2091<=SI2091;
out2092<=SI2092;
out2093<=SI2093;
out2094<=SI2094;
out2095<=SI2095;
out2096<=SI2096;
out2097<=SI2097;
out2098<=SI2098;
out2099<=SI2099;
out2100<=SI2100;
out2101<=SI2101;
out2102<=SI2102;
out2103<=SI2103;
out2104<=SI2104;
out2105<=SI2105;
out2106<=SI2106;
out2107<=SI2107;
out2108<=SI2108;
out2109<=SI2109;
out2110<=SI2110;
out2111<=SI2111;
out2112<=SI2112;
out2113<=SI2113;
out2114<=SI2114;
out2115<=SI2115;
out2116<=SI2116;
out2117<=SI2117;
out2118<=SI2118;
out2119<=SI2119;
out2120<=SI2120;
out2121<=SI2121;
out2122<=SI2122;
out2123<=SI2123;
out2124<=SI2124;
out2125<=SI2125;
out2126<=SI2126;
out2127<=SI2127;
out2128<=SI2128;
out2129<=SI2129;
out2130<=SI2130;
out2131<=SI2131;
out2132<=SI2132;
out2133<=SI2133;
out2134<=SI2134;
out2135<=SI2135;
out2136<=SI2136;
out2137<=SI2137;
out2138<=SI2138;
out2139<=SI2139;
out2140<=SI2140;
out2141<=SI2141;
out2142<=SI2142;
out2143<=SI2143;
out2144<=SI2144;
out2145<=SI2145;
out2146<=SI2146;
out2147<=SI2147;
out2148<=SI2148;
out2149<=SI2149;
out2150<=SI2150;
out2151<=SI2151;
out2152<=SI2152;
out2153<=SI2153;
out2154<=SI2154;
out2155<=SI2155;
out2156<=SI2156;
out2157<=SI2157;
out2158<=SI2158;
out2159<=SI2159;
out2160<=SI2160;
out2161<=SI2161;
out2162<=SI2162;
out2163<=SI2163;
out2164<=SI2164;
out2165<=SI2165;
out2166<=SI2166;
out2167<=SI2167;
out2168<=SI2168;
out2169<=SI2169;
out2170<=SI2170;
out2171<=SI2171;
out2172<=SI2172;
out2173<=SI2173;
out2174<=SI2174;
out2175<=SI2175;
out2176<=SI2176;
out2177<=SI2177;
out2178<=SI2178;
out2179<=SI2179;
out2180<=SI2180;
out2181<=SI2181;
out2182<=SI2182;
out2183<=SI2183;
out2184<=SI2184;
out2185<=SI2185;
out2186<=SI2186;
out2187<=SI2187;
out2188<=SI2188;
out2189<=SI2189;
out2190<=SI2190;
out2191<=SI2191;
out2192<=SI2192;
out2193<=SI2193;
out2194<=SI2194;
out2195<=SI2195;
out2196<=SI2196;
out2197<=SI2197;
out2198<=SI2198;
out2199<=SI2199;
out2200<=SI2200;
out2201<=SI2201;
out2202<=SI2202;
out2203<=SI2203;
out2204<=SI2204;
out2205<=SI2205;
out2206<=SI2206;
out2207<=SI2207;
out2208<=SI2208;
out2209<=SI2209;
out2210<=SI2210;
out2211<=SI2211;
out2212<=SI2212;
out2213<=SI2213;
out2214<=SI2214;
out2215<=SI2215;
out2216<=SI2216;
out2217<=SI2217;
out2218<=SI2218;
out2219<=SI2219;
out2220<=SI2220;
out2221<=SI2221;
out2222<=SI2222;
out2223<=SI2223;
out2224<=SI2224;
out2225<=SI2225;
out2226<=SI2226;
out2227<=SI2227;
out2228<=SI2228;
out2229<=SI2229;
out2230<=SI2230;
out2231<=SI2231;
out2232<=SI2232;
out2233<=SI2233;
out2234<=SI2234;
out2235<=SI2235;
out2236<=SI2236;
out2237<=SI2237;
out2238<=SI2238;
out2239<=SI2239;
out2240<=SI2240;
out2241<=SI2241;
out2242<=SI2242;
out2243<=SI2243;
out2244<=SI2244;
out2245<=SI2245;
out2246<=SI2246;
out2247<=SI2247;
out2248<=SI2248;
out2249<=SI2249;
out2250<=SI2250;
out2251<=SI2251;
out2252<=SI2252;
out2253<=SI2253;
out2254<=SI2254;
out2255<=SI2255;
out2256<=SI2256;
out2257<=SI2257;
out2258<=SI2258;
out2259<=SI2259;
out2260<=SI2260;
out2261<=SI2261;
out2262<=SI2262;
out2263<=SI2263;
out2264<=SI2264;
out2265<=SI2265;
out2266<=SI2266;
out2267<=SI2267;
out2268<=SI2268;
out2269<=SI2269;
out2270<=SI2270;
out2271<=SI2271;
out2272<=SI2272;
out2273<=SI2273;
out2274<=SI2274;
out2275<=SI2275;
out2276<=SI2276;
out2277<=SI2277;
out2278<=SI2278;
out2279<=SI2279;
out2280<=SI2280;
out2281<=SI2281;
out2282<=SI2282;
out2283<=SI2283;
out2284<=SI2284;
out2285<=SI2285;
out2286<=SI2286;
out2287<=SI2287;
out2288<=SI2288;
out2289<=SI2289;
out2290<=SI2290;
out2291<=SI2291;
out2292<=SI2292;
out2293<=SI2293;
out2294<=SI2294;
out2295<=SI2295;
out2296<=SI2296;
out2297<=SI2297;
out2298<=SI2298;
out2299<=SI2299;
out2300<=SI2300;
out2301<=SI2301;
out2302<=SI2302;
out2303<=SI2303;
out2304<=SI2304;
END;